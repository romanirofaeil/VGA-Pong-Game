library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity Game is
    Port(
        clk, reset, left_player, right_player : in std_logic;
        H_sync, V_sync : out std_logic;
        R_out, G_out, B_out : out std_logic_vector(3 downto 0)
        );
end Game;

architecture Behavioral of Game is

signal H_counter, V_counter, clk_counter : integer := 0;
signal image_counter : integer range 0 to 9999 := 0;
signal V_ball_move : integer range -2250 to 2250 := 0;
signal H_ball_move : integer range -3050 to 3050 := 0;
signal left_move, right_move : integer range -170 to 170 := 0;
signal sub_clk : std_logic := '0';
signal ball_down, ball_right : boolean := true;
signal end_game : boolean := false;

type data is array (0 to 9999) of STD_LOGIC_VECTOR(3 downto 0);
signal image_R: data:=("0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0001","0001","0010","0010","0001","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","0111","1001","1010","1010","1001","1001","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1001","1000","0100","0011","0100","0100","0100","0101","0100","0101","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","1001","1000","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1000","1000","0010","0001","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0001","0001","0001","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0001","0001","0001","0001","0001","0010","0101","1010","0011","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0011","1001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0101","1000","0010","0000","0000","0000","0000","0000","0000","0001","0001","0000","0000","0000","0100","0111","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1000","0101","0000","0000","0000","0000","0000","0000","0001","0001","0000","0000","0000","0110","0101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","0111","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0110","0101","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0100","0101","0110","0110","0101","0100","0011","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0100","0100","0010","0010","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0010","0011","0010","0001","0000","0000","0000","0000","0001","0001","0010","0010","0001","0001","0000","0000","0000","0000","0000","0001","0001","0001","0010","0001","0001","0001","0010","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0010","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0110","0101","0000","0001","0000","0000","0000","0000","0000","0001","0011","0110","1001","1101","1111","1111","1111","1011","0111","0100","0010","0001","0001","0000","0000","0000","0000","0000","0000","0000","0001","0011","0110","1000","1000","0110","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0011","0110","0111","0110","0011","0001","0000","0000","0001","0010","0100","0110","0101","0100","0011","0001","0000","0000","0000","0000","0001","0010","0100","0100","0100","0100","0101","0100","0101","0100","0100","0011","0001","0001","0000","0000","0000","0000","0010","1000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0110","0101","0000","0000","0000","0000","0000","0001","0001","0100","1000","1101","1111","1111","1100","1011","1100","1111","1111","1010","0101","0010","0001","0000","0000","0000","0000","0000","0001","0000","0010","0110","1101","1111","1111","1101","0110","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","1000","1101","1111","1101","1000","0011","0001","0001","0010","0110","1010","1100","1011","1001","0101","0011","0001","0000","0000","0000","0011","1001","1110","1110","1110","1110","1110","1110","1110","1110","1110","1100","0110","0010","0001","0000","0000","0000","0011","1000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0110","0101","0000","0000","0000","0000","0000","0010","0100","1001","1111","1101","1000","0111","0110","0110","0110","0111","1011","1111","1011","0101","0010","0001","0000","0000","0000","0000","0000","0001","0100","1100","1110","1001","1000","1111","1011","0011","0001","0000","0000","0000","0000","0000","0000","0000","0001","0001","0101","1110","1110","1100","1101","1111","0110","0010","0010","0100","1010","1111","1110","1110","1111","1000","0011","0001","0000","0000","0001","1001","1110","1000","1000","0111","1000","1000","0111","1000","1000","1000","1010","1110","0100","0001","0000","0000","0000","0011","1000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0110","0101","0000","0000","0000","0000","0001","0011","1000","1111","1100","0110","0100","0100","0101","0101","0100","0100","0110","1010","1111","1011","0101","0010","0000","0000","0000","0000","0001","0010","0110","1111","1001","0100","0100","1001","1111","0101","0010","0001","0000","0000","0000","0000","0000","0000","0001","0010","0111","1111","1000","0101","0111","1111","1001","0011","0010","0110","1110","1011","0110","0111","1101","1010","0011","0001","0001","0001","0010","1110","0111","0010","0000","0001","0001","0001","0010","0001","0010","0010","0011","1101","0101","0001","0000","0000","0000","0011","1000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0110","0101","0000","0000","0000","0000","0010","0110","1111","1100","0111","0100","0101","0110","1000","1000","0111","0101","0100","0101","1010","1111","1001","0011","0001","0000","0000","0000","0001","0100","1010","1111","0110","0010","0010","0110","1111","1000","0011","0001","0000","0000","0000","0000","0000","0001","0001","0011","1000","1110","0101","0011","0100","1100","1100","0100","0011","1000","1111","1000","0100","0100","1010","1100","0101","0001","0000","0001","0011","1111","0101","0001","0000","0010","0010","0010","0010","0010","0011","0011","0100","1110","0101","0001","0000","0000","0000","0011","1000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0110","0101","0000","0000","0000","0001","0011","1001","1111","0111","0100","0101","1000","1110","1111","1111","1111","1010","0101","0011","0100","1010","1111","0101","0010","0001","0000","0001","0010","0101","1110","1010","0100","0010","0001","0101","1100","1011","0100","0001","0000","0000","0000","0000","0000","0000","0001","0100","1011","1100","0101","0010","0010","1000","1111","0110","0101","1011","1111","0101","0011","0011","1000","1110","0110","0001","0000","0000","0011","1110","0100","0010","0001","0111","1011","1011","1011","1100","1100","1100","1101","1101","0011","0001","0000","0000","0000","0010","1000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0110","0101","0000","0000","0001","0001","0100","1101","1011","0100","0011","1000","1111","1110","1000","1000","1100","1111","1000","0010","0011","0110","1111","0111","0010","0001","0001","0001","0010","0111","1111","0111","0011","0001","0010","0011","1000","1111","0110","0010","0001","0000","0000","0000","0000","0000","0010","0100","1101","1010","0011","0001","0010","0110","1111","1001","0111","1111","1010","0011","0001","0010","0110","1111","0110","0010","0000","0000","0011","1110","0100","0001","0011","1101","1111","1110","1101","1110","1101","1101","1100","0101","0010","0001","0000","0000","0000","0010","1000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0110","0101","0000","0000","0001","0010","0101","1111","1000","0010","0011","1100","1111","0110","0100","0011","0101","1101","1101","0110","0100","0110","1110","1000","0011","0001","0001","0001","0100","1011","1101","0100","0010","0011","0011","0011","0110","1111","1001","0011","0001","0000","0000","0000","0000","0001","0010","0110","1111","1000","0011","0001","0001","0101","1101","1101","1001","1111","0111","0010","0001","0001","0100","1111","1001","0010","0001","0001","0010","1111","0100","0001","0010","1110","0110","0010","0010","0010","0010","0010","0010","0001","0001","0000","0000","0000","0000","0010","1001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0110","0101","0000","0000","0000","0010","0101","1111","1000","0010","0011","1110","1010","0100","0010","0001","0010","1000","1111","1000","0111","1001","1111","0111","0010","0001","0001","0010","0101","1111","1001","0100","0011","0110","0110","0100","0101","1011","1101","0101","0010","0000","0000","0000","0000","0000","0010","1000","1111","0110","0010","0001","0001","0011","1001","1111","1100","1110","0100","0001","0000","0001","0011","1110","1010","0011","0001","0001","0011","1110","0101","0001","0010","1110","0100","0001","0001","0001","0010","0001","0001","0000","0000","0000","0000","0000","0000","0011","1001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0101","0101","0000","0000","0000","0010","0101","1111","0111","0010","0100","1110","1010","0011","0001","0001","0010","0110","1111","1111","1110","1111","1100","0100","0010","0000","0001","0011","1001","1111","0111","0011","0110","1111","1110","0110","0101","1000","1111","0111","0010","0000","0000","0000","0000","0000","0010","1001","1110","0100","0001","0001","0001","0010","0110","1111","1111","1001","0011","0001","0001","0000","0010","1011","1101","0100","0010","0001","0011","1110","0101","0010","0010","1110","0110","0011","0011","0011","0010","0010","0001","0000","0000","0000","0000","0000","0000","0011","1001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0101","0101","0000","0000","0000","0010","0101","1111","0111","0010","0100","1110","1001","0010","0001","0010","0101","0110","1001","1100","1101","1011","0111","0011","0001","0001","0001","0101","1110","1011","0101","0101","1001","1111","1111","1001","0101","0110","1101","1011","0100","0001","0000","0000","0000","0001","0011","1011","1100","0011","0001","0001","0010","0010","0100","1001","1100","0101","0010","0001","0001","0001","0010","1000","1110","0110","0010","0010","0011","1110","0100","0001","0010","1100","1110","1101","1100","1100","1100","1000","0010","0000","0000","0000","0000","0000","0000","0010","1001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0101","0101","0000","0000","0000","0010","0110","1111","0110","0011","0100","1110","1001","0100","0100","0111","1001","1010","1011","1010","1010","1001","0110","0010","0010","0001","0010","0111","1111","0111","0100","0110","1101","1101","1101","1110","0110","0101","1001","1110","0101","0001","0000","0000","0000","0001","0100","1101","1010","0011","0010","0011","0011","0010","0010","0100","0100","0001","0001","0011","0011","0010","0011","0111","1111","0110","0010","0010","0011","1110","0100","0001","0000","0101","1001","1010","1011","1011","1100","1111","0111","0001","0000","0000","0000","0000","0000","0010","1001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0101","0110","0000","0000","0000","0010","0110","1111","0110","0011","0100","1110","1010","0100","1001","1111","1111","1111","1111","1111","1111","1111","1010","0100","0010","0010","0100","1011","1101","0101","0011","1000","1111","1010","1010","1111","1000","0100","0110","1111","1000","0010","0001","0000","0001","0010","0101","1111","1001","0011","0011","0111","1010","0100","0010","0010","0001","0000","0001","0101","1010","0101","0011","0110","1111","0111","0011","0010","0011","1110","0100","0000","0001","0010","0011","0011","0011","0011","0011","1001","1100","0001","0000","0000","0000","0000","0000","0011","1001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0101","0110","0000","0000","0000","0011","0110","1111","0110","0010","0100","1110","1001","0110","1101","1100","1000","1000","0111","1000","1000","1011","1111","0110","0011","0010","0101","1111","1010","0011","0011","1011","1110","1001","1001","1111","1001","0011","0100","1100","1100","0100","0010","0001","0001","0011","0111","1111","0111","0010","0100","1101","1111","1000","0011","0001","0001","0001","0100","1011","1111","1000","0101","0101","1101","1010","0100","0010","0011","1110","0100","0001","0001","0010","0011","0011","0011","0100","0011","1001","1100","0001","0001","0001","0000","0000","0000","0011","1010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0101","0110","0000","0000","0001","0010","0111","1111","0110","0010","0101","1111","1010","0110","1111","1010","0111","0110","0101","0100","0100","0111","1111","1000","0011","0100","1000","1111","0110","0010","0011","1011","1111","1111","1111","1111","1010","0011","0011","1000","1111","0110","0011","0001","0001","0100","1000","1111","0101","0011","0101","1111","1101","1100","0100","0001","0001","0010","0110","1111","1110","1011","0101","0101","1011","1101","0101","0001","0011","1110","0100","0001","0001","0100","0111","0111","0111","0110","0111","1110","1001","0001","0000","0000","0000","0000","0000","0011","1010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0101","0110","0000","0000","0001","0010","0110","1111","0110","0011","0101","1111","1010","0110","1100","1110","1010","1010","0111","0011","0011","0110","1101","1000","0100","0101","1101","1011","0100","0010","0010","0110","1010","1011","1011","1010","0110","0001","0010","0101","1110","1001","0011","0001","0001","0100","1011","1100","0100","0011","0111","1111","1011","1111","0110","0010","0001","0011","1000","1111","1100","1101","0101","0100","1000","1111","0101","0010","0011","1110","0100","0001","0010","1011","1110","1110","1110","1110","1101","1101","0100","0001","0000","0000","0000","0000","0000","0010","1010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0101","0110","0000","0001","0000","0010","0101","1111","0110","0011","0100","1111","1001","0101","1000","1110","1111","1111","1110","0100","0011","0101","1111","1000","0100","0111","1111","1000","0011","0010","0010","0100","0101","0101","0101","0101","0011","0010","0010","0100","1011","1101","0101","0001","0001","0101","1101","1010","0100","0100","1010","1110","1001","1111","1000","0011","0011","0100","1101","1101","1010","1111","0101","0100","0111","1111","0111","0010","0011","1110","0101","0001","0010","1111","0110","0100","0100","0100","0100","0011","0010","0000","0000","0000","0000","0000","0000","0010","1010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0101","0110","0000","0000","0000","0001","0101","1111","1000","0011","0100","1100","1101","0111","0110","1000","1010","1100","1111","0101","0011","0111","1111","1000","0101","1011","1110","0100","0010","0011","0101","0110","0110","0111","0110","0110","0101","0100","0011","0011","0111","1111","0111","0010","0010","0110","1111","1000","0100","0100","1100","1011","0111","1110","1011","0101","0101","1000","1111","1010","1000","1111","0110","0011","0101","1111","1000","0011","0011","1110","0100","0001","0010","1110","0100","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","1001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0101","0110","0000","0000","0000","0001","0100","1110","1010","0100","0011","1000","1111","1101","1001","1001","1011","1111","1011","0100","0011","1000","1111","1000","0111","1111","1010","0011","0011","0110","1110","1110","1110","1111","1111","1110","1101","1011","0101","0011","0101","1110","1010","0011","0010","0111","1111","0110","0011","0110","1110","1000","0101","1010","1111","1100","1010","1111","1111","0111","0111","1111","0111","0011","0100","1110","1010","0011","0100","1110","0100","0001","0010","1110","0101","0010","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0010","1001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0101","0111","0000","0000","0000","0001","0011","1010","1110","0110","0100","0101","1001","1111","1111","1111","1111","1100","0110","0011","0100","1011","1110","0111","1000","1111","0111","0010","0100","1100","1111","1101","1101","1101","1110","1110","1111","1111","1000","0100","0100","1001","1111","0101","0011","1000","1111","0101","0011","0111","1111","0110","0100","0110","1011","1111","1111","1111","1000","0100","0101","1110","1001","0100","0100","1100","1100","0100","0101","1110","0100","0001","0010","1111","1010","1000","1000","0111","0110","0110","0110","0010","0001","0000","0000","0000","0000","0010","1010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0101","0111","0000","0000","0000","0001","0010","0110","1111","1011","0110","0100","0101","0111","1001","1010","1000","0110","0100","0100","1000","1111","1001","0110","1100","1110","0101","0011","0110","1111","1010","0110","0110","0110","0110","0101","0111","1100","1101","0100","0011","0111","1111","1000","0100","1011","1110","0100","0011","1000","1111","0110","0011","0011","0101","0110","0110","0110","0100","0010","0011","1101","1011","0100","0011","1001","1111","0101","0101","1111","0100","0001","0010","1010","1111","1111","1111","1110","1111","1111","1110","1001","0010","0001","0000","0000","0000","0010","1010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0101","0110","0000","0000","0000","0000","0001","0011","1000","1111","1010","0111","0100","0100","0100","0100","0100","0100","0110","0111","1110","1100","0111","0110","1111","1011","0101","0110","1010","1110","0110","0011","0001","0001","0010","0010","0011","0111","1111","0111","0100","0110","1101","1010","0110","1101","1100","0101","0101","1011","1110","0100","0010","0001","0001","0010","0010","0001","0001","0001","0010","1011","1101","0101","0011","0111","1111","0110","0101","1110","0100","0001","0000","0001","0011","0011","0011","0100","0100","0100","0110","1110","0100","0001","0000","0000","0000","0010","1010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","0110","0000","0000","0000","0000","0000","0010","0101","1010","1111","1011","1000","0101","0101","0101","0110","0111","1010","1111","1110","0111","0100","0101","1101","1100","1000","1001","1110","1011","0011","0001","0000","0000","0000","0000","0001","0101","1110","1011","0110","0111","1110","1010","0110","1100","1100","0111","0111","1101","1100","0011","0001","0000","0000","0000","0000","0000","0000","0000","0010","1001","1111","0110","0100","0111","1111","0110","0101","1111","0101","0001","0001","0001","0001","0001","0001","0001","0001","0010","0011","1101","0100","0001","0000","0000","0000","0010","1010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","0110","0000","0000","0000","0000","0000","0001","0010","0101","1001","1111","1111","1110","1110","1101","1101","1111","1111","1100","0110","0010","0010","0011","1001","1111","1111","1111","1110","0110","0010","0001","0000","0000","0000","0000","0001","0011","1001","1111","1110","1110","1111","0111","0100","1000","1111","1110","1110","1111","0111","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","0110","1111","1101","1010","1101","1110","0100","0011","1101","1011","0110","0101","0101","0100","0100","0100","0100","0100","0100","0110","1110","0100","0001","0000","0000","0000","0010","1010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","0110","0000","0000","0000","0000","0000","0000","0001","0011","0100","0111","1010","1101","1110","1111","1110","1011","1000","0101","0010","0001","0000","0010","0101","1001","1101","1011","0111","0011","0001","0000","0000","0000","0000","0000","0001","0010","0101","1010","1110","1111","1001","0011","0010","0101","1001","1101","1100","1001","0100","0001","0000","0000","0000","0000","0000","0000","0000","0001","0001","0100","1001","1111","1111","1111","0111","0011","0010","0101","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1010","0010","0001","0000","0000","0000","0010","1010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","0111","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0100","0101","0110","0110","0110","0100","0011","0010","0001","0000","0000","0000","0001","0100","0100","0100","0010","0001","0000","0000","0000","0001","0000","0000","0000","0000","0010","0100","0110","0101","0100","0010","0001","0010","0011","0101","0101","0011","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0100","0110","0111","0110","0011","0001","0001","0001","0011","0111","0111","0111","1000","1000","1000","1000","1000","1000","0111","0011","0001","0000","0000","0000","0000","0010","1010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","0111","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0011","0100","0100","0100","0011","0010","0001","0001","0001","0000","0000","0000","0001","0010","0010","0001","0001","0000","0000","0001","0000","0000","0000","0000","0000","0000","0001","0010","0010","0010","0001","0001","0010","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0010","0010","0011","0011","0011","0010","0001","0010","0010","0011","0011","0100","0011","0100","0011","0011","0011","0010","0010","0001","0001","0000","0000","0000","0000","0000","0010","1010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","0111","0000","0000","0000","0000","0000","0000","0001","0000","0000","0001","0011","0110","1000","1001","1000","0111","0101","0011","0010","0001","0000","0000","0000","0000","0010","0011","0011","0010","0001","0001","0000","0000","0000","0000","0001","0000","0000","0001","0001","0001","0010","0010","0010","0010","0001","0001","0001","0011","0100","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0011","0010","0010","0010","0011","0101","0110","0111","0110","0111","0111","0111","0111","0110","0101","0011","0010","0010","0001","0000","0001","0000","0000","0000","0000","0010","1010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","0111","0000","0000","0000","0000","0001","0001","0000","0001","0010","0110","1100","1111","1111","1111","1111","1110","1110","1100","0111","0010","0001","0000","0000","0001","0100","1011","1101","1010","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0101","1010","1100","0111","0010","0001","0001","0101","1010","1110","1110","1111","1111","1111","1110","1110","1111","1110","1110","1101","1000","0011","0010","0011","0110","1011","1110","1111","1111","1110","1110","1111","1101","1100","1001","0110","0011","0010","0001","0000","0000","0000","0000","0000","0000","0010","1010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","0111","0000","0000","0000","0000","0000","0001","0001","0011","1001","1111","1011","0110","0100","0011","0011","0100","0110","1010","1111","1001","0010","0001","0001","0011","1011","1101","1001","1100","1100","0010","0001","0000","0000","0000","0000","0000","0000","0000","0001","0011","1110","1100","1011","1111","0110","0010","0011","1010","1111","1100","1100","1100","1100","1100","1100","1100","1100","1011","1100","1101","1111","0101","0011","0101","1101","1111","1101","1100","1100","1100","1101","1100","1110","1111","1111","1110","1000","0101","0010","0001","0000","0000","0000","0000","0000","0010","1010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","0111","0000","0000","0000","0000","0001","0001","0010","1000","1111","0111","0011","0011","0010","0001","0001","0010","0010","0011","0111","1111","1001","0010","0010","0011","1110","0110","0011","0101","1110","0101","0001","0000","0000","0000","0000","0000","0000","0000","0001","1000","1101","0100","0011","1001","1100","0011","0101","1111","1011","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","1000","1111","1000","0011","0110","1111","1001","0110","0110","0111","0110","0110","0111","0111","0111","1000","1101","1111","1010","0101","0001","0000","0000","0000","0000","0000","0010","1010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","0111","0000","0000","0000","0000","0001","0010","0111","1110","0110","0010","0010","0011","0100","0101","0100","0100","0011","0001","0001","0110","1110","1000","0010","0011","1101","0101","0010","0010","1001","1001","0010","0001","0000","0000","0000","0000","0001","0001","0010","1100","0111","0010","0010","1000","1101","0100","0111","1111","0111","0011","0011","0101","0111","1000","1000","1000","1000","1000","0111","1001","1111","1000","0011","0111","1111","0110","0100","0100","0101","0110","0111","0111","0110","0101","0101","0110","1010","1111","1001","0011","0001","0000","0000","0000","0000","0010","1010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","0111","0000","0000","0000","0000","0001","0100","1110","1000","0011","0001","0010","0111","1110","1111","1111","1110","1000","0001","0001","0010","1000","1111","0101","0011","1100","0110","0010","0010","0101","1101","0011","0001","0000","0000","0000","0001","0000","0001","0100","1110","0100","0001","0010","1100","1001","0100","1000","1111","0110","0010","0011","0111","1010","1010","1010","1011","1010","1010","1010","1011","1111","0101","0011","0110","1111","0110","0011","0100","1000","1011","1011","1011","1001","0111","0101","0100","0110","1010","1111","0101","0010","0000","0000","0000","0000","0010","1010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","1000","0000","0000","0000","0000","0010","1000","1101","0011","0010","0010","1000","1110","1011","0111","0111","1011","1111","1010","0010","0010","0011","1101","1011","0011","1000","1011","0010","0001","0011","1110","0101","0010","0000","0000","0000","0000","0000","0001","1000","1011","0010","0010","0100","1110","0101","0100","1000","1110","0110","0011","0100","1101","1111","1111","1111","1111","1111","1111","1111","1111","1001","0011","0010","0110","1111","0110","0011","0110","1111","1111","1111","1111","1111","1111","1001","0100","0100","0110","1111","1001","0011","0000","0000","0000","0000","0010","1010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","1000","0001","0000","0000","0000","0010","1100","0111","0010","0010","0111","1110","0111","0011","0010","0010","0011","0110","1110","1000","0010","0010","0111","1110","0011","0101","1110","0101","0001","0001","1010","1001","0010","0000","0000","0000","0000","0000","0010","1101","0110","0010","0010","1000","1100","0011","0100","1000","1110","0110","0011","0110","1111","1001","0101","0101","0101","0101","0101","0101","0101","0011","0001","0010","0101","1111","0101","0100","0110","1111","1001","0111","0110","0111","1011","1111","0111","0011","0101","1001","1110","0100","0001","0000","0000","0000","0001","1010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","1000","0001","0000","0000","0001","0010","1101","0100","0010","0011","1100","1000","0001","0001","0001","0001","0001","0010","1000","1101","0001","0001","0100","1110","0100","0010","1101","1000","0001","0001","0110","1101","0011","0001","0001","0000","0000","0000","0101","1110","0010","0001","0011","1101","0111","0010","0100","1000","1110","0110","0100","0110","1111","0110","0010","0001","0001","0001","0010","0001","0001","0000","0000","0001","0110","1111","0110","0011","0110","1111","0111","0100","0010","0010","0110","1110","1001","0100","0011","0110","1111","0110","0001","0000","0000","0000","0001","1010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","1000","0001","0000","0000","0001","0011","1101","0100","0010","0011","1101","0100","0001","0000","0000","0000","0000","0001","0101","1101","0001","0001","0011","1110","0011","0010","1001","1101","0010","0001","0011","1101","0110","0010","0001","0000","0000","0001","1010","1011","0001","0001","0101","1110","0011","0010","0011","1000","1110","0110","0100","0111","1111","0110","0010","0001","0001","0001","0001","0001","0001","0000","0000","0001","0110","1111","0110","0011","0111","1111","0111","0011","0001","0001","0100","1100","1011","0100","0011","0101","1111","0110","0010","0000","0000","0000","0001","1010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","1000","0001","0000","0000","0000","0011","1110","0011","0010","0011","1110","0100","0000","0000","0000","0001","0000","0001","0101","1110","0001","0001","0011","1101","0011","0010","0100","1111","0100","0010","0010","1001","1001","0010","0001","0001","0001","0011","1110","0101","0010","0010","1010","1011","0010","0001","0011","1000","1110","0110","0011","0111","1111","0111","0011","0010","0011","0011","0011","0010","0001","0000","0000","0001","0110","1111","0110","0011","0111","1110","0111","0011","0010","0010","0100","1011","1011","0101","0011","0101","1111","0111","0010","0000","0000","0000","0001","1010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","1000","0001","0000","0000","0001","0011","1110","0011","0001","0011","1110","0011","0001","0000","0000","0000","0000","0000","0101","1110","0001","0001","0100","1101","0011","0010","0011","1011","1000","0010","0010","0101","1101","0100","0001","0000","0001","0111","1101","0011","0010","0011","1110","0110","0010","0001","0011","1000","1110","0110","0011","0110","1111","1001","1000","1000","0111","0111","0111","0101","0011","0001","0001","0010","0110","1111","0110","0100","0111","1111","0111","0100","0011","0011","0110","1111","1000","0100","0011","0110","1111","0110","0010","0000","0000","0000","0001","1010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","1000","0001","0000","0000","0001","0011","1101","0011","0001","0010","1110","0011","0001","0000","0000","0000","0000","0001","0101","1110","0001","0001","0100","1110","0100","0010","0010","0111","1101","0011","0001","0010","1110","0111","0001","0001","0011","1011","1000","0010","0010","0111","1101","0011","0001","0001","0011","1000","1110","0101","0010","0100","1101","1111","1111","1111","1111","1111","1111","1101","0101","0010","0001","0001","0110","1111","0110","0100","0110","1111","1010","1000","1000","1001","1110","1101","0101","0011","0100","1001","1111","0101","0001","0000","0000","0000","0001","1001","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","1000","0001","0000","0000","0001","0011","1101","0011","0001","0010","1101","0011","0001","0000","0000","0000","0000","0001","0101","1110","0001","0001","0011","1110","0100","0010","0010","0100","1111","0101","0001","0001","1010","1011","0010","0010","0100","1111","0100","0010","0011","1010","1000","0010","0001","0001","0011","1000","1110","0101","0010","0010","0110","1001","1001","1010","1010","1010","1010","1111","1000","0011","0001","0010","0110","1111","0110","0011","0101","1110","1111","1111","1111","1111","1100","0111","0011","0010","0110","1100","1011","0100","0001","0000","0000","0000","0001","1001","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","1000","0001","0000","0000","0001","0011","1101","0010","0001","0010","1101","0011","0001","0000","0000","0000","0000","0001","0101","1110","0000","0000","0011","1110","0011","0001","0001","0010","1011","1010","0001","0001","0101","1110","0011","0010","1001","1101","0011","0001","0100","1110","0100","0001","0000","0001","0011","1000","1110","0101","0001","0001","0011","0101","0110","0101","0101","0101","0111","1011","1100","0011","0001","0001","0110","1111","0101","0011","0011","0110","1000","1000","1000","0111","0110","0011","0010","0011","1000","1111","0111","0010","0001","0000","0000","0000","0001","1001","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1000","0001","0000","0000","0001","0011","1110","0010","0001","0010","1101","0011","0000","0000","0000","0000","0000","0001","0110","1110","0000","0000","0011","1101","0100","0001","0001","0001","0110","1110","0010","0001","0011","1101","0111","0100","1101","1000","0010","0010","1000","1100","0010","0001","0000","0001","0011","1001","1110","0110","0010","0010","0101","0110","0110","0110","0110","0101","0110","1101","1011","0011","0001","0001","0110","1111","0110","0010","0010","0011","0100","0101","0101","0101","0100","0011","0010","0110","1110","1100","0101","0010","0001","0000","0000","0000","0001","1001","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1000","0001","0000","0000","0001","0100","1110","0010","0001","0011","1101","0011","0000","0000","0000","0000","0000","0001","0110","1110","0001","0000","0010","1110","0100","0001","0000","0001","0011","1110","0100","0001","0011","1001","1100","0110","1110","0100","0001","0010","1100","0111","0001","0000","0000","0001","0011","1001","1111","0110","0011","0100","1010","1100","1100","1100","1011","1011","1100","1111","1000","0011","0001","0001","0110","1111","0101","0010","0011","0100","0110","0111","0110","0110","0100","0100","0011","0111","1111","1000","0011","0010","0001","0000","0000","0000","0001","1001","0010","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0011","1000","0001","0000","0000","0001","0100","1110","0010","0001","0011","1110","0011","0000","0000","0000","0000","0000","0001","0110","1110","0010","0001","0010","1101","0100","0001","0000","0001","0010","1010","1010","0010","0010","0101","1111","1100","1011","0010","0001","0100","1110","0100","0001","0000","0000","0001","0011","1001","1110","0110","0011","0110","1111","1111","1111","1111","1111","1111","1110","1011","0100","0010","0001","0001","0110","1111","0101","0010","0100","1000","1100","1101","1100","1100","1010","0101","0011","0101","1101","1100","0011","0010","0001","0000","0000","0000","0001","1001","0010","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0011","1000","0001","0000","0000","0001","0100","1110","0010","0001","0011","1101","0011","0001","0000","0000","0000","0000","0001","0110","1110","0010","0001","0011","1101","0100","0001","0000","0001","0001","0100","1110","0011","0001","0010","1100","1111","0101","0010","0010","1000","1011","0010","0001","0000","0000","0001","0011","1000","1110","0101","0100","0111","1111","1000","0110","0101","0110","0101","0110","0100","0001","0000","0000","0010","0110","1111","0101","0011","0110","1111","1111","1111","1111","1111","1111","1000","0100","0011","1000","1111","0110","0010","0001","0000","0000","0000","0001","1001","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1000","0001","0000","0000","0001","0100","1110","0011","0001","0011","1110","0100","0001","0000","0000","0000","0001","0010","0111","1110","0001","0001","0011","1110","0011","0001","0000","0000","0001","0011","1101","0110","0001","0001","0101","0111","0010","0001","0011","1100","0110","0010","0001","0000","0000","0001","0011","1000","1110","0101","0100","0111","1111","0110","0011","0010","0010","0010","0010","0001","0000","0000","0000","0010","0111","1111","0101","0011","0110","1111","1000","0110","0110","0110","1100","1110","0100","0011","0110","1110","0110","0010","0001","0000","0000","0000","0001","1001","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1000","0001","0000","0001","0001","0011","1110","0011","0001","0010","1100","1001","0010","0001","0000","0001","0010","0100","1101","1001","0001","0001","0101","1110","0011","0001","0000","0000","0000","0001","1010","1011","0001","0001","0001","0001","0001","0001","0101","1110","0010","0001","0001","0000","0000","0001","0011","1000","1101","0110","0100","0111","1111","0110","0010","0001","0001","0001","0001","0001","0000","0000","0000","0010","0111","1111","0101","0011","0110","1111","0111","0011","0011","0011","0111","1111","0110","0011","0101","1101","0111","0011","0001","0000","0000","0000","0001","1001","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1001","0001","0000","0000","0001","0011","1101","0110","0001","0001","1000","1111","0110","0010","0010","0010","0100","1010","1110","0100","0001","0001","0111","1101","0010","0001","0000","0000","0000","0001","0110","1110","0100","0001","0000","0000","0000","0001","1010","1010","0001","0001","0001","0000","0000","0001","0011","1001","1110","0101","0100","0111","1111","0110","0010","0010","0001","0001","0001","0010","0001","0001","0001","0010","0111","1111","0101","0011","0110","1110","0110","0011","0001","0001","0110","1111","0111","0011","0101","1101","1000","0011","0001","0000","0000","0000","0001","1001","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1001","0001","0000","0000","0000","0001","1001","1010","0011","0010","0011","1001","1110","1011","1001","1010","1101","1110","0110","0010","0010","0010","1100","1001","0001","0001","0000","0000","0000","0001","0011","1101","0110","0010","0001","0000","0001","0011","1110","0110","0001","0000","0000","0000","0000","0001","0100","1000","1110","0101","0100","0110","1111","1000","0111","0111","0111","0110","0111","0110","0101","0011","0001","0010","0111","1111","0101","0011","0110","1111","0111","0011","0001","0001","0101","1111","0111","0100","0110","1110","1001","0011","0001","0000","0000","0000","0001","1001","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1001","0001","0000","0000","0000","0001","0100","1110","0111","0010","0010","0010","1000","1011","1110","1101","1010","0100","0010","0010","0011","1001","1101","0011","0001","0000","0000","0000","0000","0001","0010","1001","1011","0011","0001","0001","0001","0111","1101","0011","0001","0000","0000","0000","0000","0001","0011","1001","1110","0101","0010","0101","1100","1111","1111","1111","1111","1111","1111","1111","1111","1000","0011","0011","0111","1111","0100","0011","0111","1111","0110","0011","0001","0001","0101","1111","0111","0100","0101","1101","1001","0011","0001","0000","0000","0000","0001","1001","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1001","0001","0000","0000","0000","0000","0010","1000","1111","0111","0010","0010","0001","0010","0011","0010","0001","0001","0010","0011","1000","1111","0110","0001","0001","0000","0000","0000","0000","0000","0001","0100","1110","0100","0001","0001","0010","1011","1000","0001","0000","0000","0000","0000","0000","0001","0011","1001","1101","0110","0010","0011","0110","1000","1001","1010","1011","1010","1011","1011","1101","1111","0101","0011","0111","1111","0101","0011","0111","1111","0110","0011","0001","0001","0101","1110","1000","0100","0101","1100","1001","0011","0001","0000","0000","0000","0001","1001","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1001","0001","0000","0000","0000","0000","0001","0011","1000","1110","1000","0011","0010","0001","0001","0001","0001","0001","0100","1001","1110","1000","0001","0001","0000","0000","0000","0000","0000","0001","0001","0010","1100","1000","0010","0010","0101","1110","0100","0001","0000","0000","0000","0000","0000","0001","0011","1000","1110","0110","0100","0011","0100","0110","0110","0110","0110","0110","0110","0110","1000","1111","0110","0011","1000","1111","0110","0100","0111","1111","0110","0010","0001","0001","0101","1110","0111","0101","0101","1100","1010","0011","0001","0001","0000","0000","0001","1001","0100","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1001","0001","0000","0000","0000","0000","0001","0001","0011","0111","1111","1100","0111","0101","0100","0100","0101","0111","1100","1111","1000","0010","0001","0001","0000","0000","0000","0000","0000","0000","0001","0001","1000","1110","0110","0110","1011","1100","0010","0001","0000","0000","0000","0000","0000","0001","0010","0111","1111","1001","0111","0111","0111","0111","0111","1000","1000","0111","0111","0111","1000","1111","0110","0011","0111","1111","1000","1000","1001","1111","0101","0001","0001","0001","0100","1110","1010","1000","1000","1110","1001","0011","0001","0000","0000","0000","0001","1000","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","1001","0001","0000","0000","0000","0000","0001","0001","0001","0010","0110","1101","1111","1110","1101","1110","1110","1111","1100","0101","0010","0010","0000","0000","0000","0000","0000","0000","0001","0000","0000","0001","0011","1100","1111","1111","1111","0110","0010","0001","0000","0000","0000","0000","0000","0001","0010","0100","1101","1111","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1111","1101","0100","0010","0101","1111","1110","1101","1111","1100","0011","0001","0000","0001","0011","1011","1111","1101","1101","1111","0110","0010","0001","0000","0000","0000","0001","1000","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1001","0001","0000","0000","0000","0000","0000","0000","0001","0001","0001","0010","0101","0110","0111","0111","0111","0100","0010","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0010","0101","0101","0011","0010","0001","0001","0000","0000","0000","0000","0000","0001","0001","0010","0101","1010","1100","1101","1101","1101","1101","1101","1101","1101","1101","1100","1011","0111","0010","0001","0011","0111","1100","1101","1011","0110","0010","0000","0000","0001","0010","0110","1011","1110","1101","1001","0100","0001","0001","0000","0000","0000","0001","1000","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1001","0001","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0010","0011","0101","0101","0110","0110","0110","0101","0101","0110","0110","0110","0101","0011","0000","0000","0001","0011","0101","0101","0100","0010","0001","0001","0000","0001","0001","0010","0101","0101","0101","0100","0001","0000","0000","0000","0000","0000","0001","1000","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1000","0100","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0000","0000","0000","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0001","1001","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0101","1001","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","1010","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0111","1001","0110","0011","0010","0001","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0001","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0110","0111","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0101","0111","1000","1000","1000","0011","0000","0000","0000","0100","0111","0101","0010","0000","0000","0001","0110","0111","1001","1001","1001","1000","1000","1000","1000","1001","1000","0101","0000","0000","0000","0001","0100","0111","0110","0010","0000","0000","0000","0000","0100","0101","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0000","0000","0000","0000","0010","0011","0010","0000","0000","0000","0000","0000","0000","0010","0011","0100","0111","1000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0001","0001","0010","0110","0110","0001","0000","0010","1010","0110","1010","0100","0000","0000","0010","1001","0101","0101","0100","0101","0101","0101","0100","0100","0101","0110","1001","0010","0000","0000","0100","1010","0111","1000","1010","0010","0000","0000","0011","1011","1001","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","0100","0000","0000","0010","1010","1011","1010","0100","0000","0000","0000","0000","0011","1010","1100","1011","0111","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1000","0000","0000","0011","0111","0001","0101","0111","0000","0000","0011","1000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0001","1000","0001","0000","0000","0111","0101","0001","0001","1000","0100","0000","0000","0101","0110","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0001","0001","0010","0010","0010","0010","0001","0010","0001","0010","0100","1000","0001","0000","0100","0111","0010","0110","1000","0000","0000","0000","0000","0110","0110","0010","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1000","0000","0000","0011","0111","0000","0100","0111","0000","0000","0010","0111","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1000","0010","0000","0000","1000","0011","0000","0000","0111","0100","0000","0000","0101","0101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1000","0000","0000","0101","0101","0000","0010","1001","0001","0000","0000","0000","0110","0100","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","1000","0000","0000","0100","0111","0000","0010","1001","0001","0000","0100","0110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1000","0010","0000","0000","1000","0011","0000","0000","0111","0100","0000","0000","0101","0101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","1001","0000","0000","0101","0100","0000","0010","1001","0001","0000","0000","0000","0110","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1000","0000","0000","0011","0110","0000","0001","1000","1000","1000","1001","0100","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1000","0010","0000","0000","1000","0100","0000","0000","0110","0101","0000","0000","0101","0101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","1001","0001","0001","0110","0100","0000","0010","1001","0001","0000","0000","0000","0110","0100","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1000","0000","0000","0100","0110","0000","0000","0010","0101","0110","0100","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1000","0010","0000","0000","1001","0011","0000","0000","0110","0101","0000","0000","0101","0101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1001","1000","0111","1001","0001","0000","0010","1010","0001","0000","0000","0000","0110","0100","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","0111","0000","0000","0011","0110","0000","0000","0000","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1000","0010","0000","0000","1001","0100","0000","0000","0101","0110","0001","0000","0110","0100","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1000","1000","0011","0000","0000","0010","1010","0001","0000","0000","0000","0110","0100","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1000","0000","0000","0100","0110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1000","0010","0000","0000","1001","0011","0000","0000","0010","1001","0111","0110","1001","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0000","0000","0010","1010","0001","0000","0000","0000","0110","0100","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1010","0100","0011","1000","0100","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1000","0001","0000","0000","1000","0100","0000","0000","0001","0100","0111","1000","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0010","1010","0001","0000","0000","0000","0111","0100","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0110","1010","1010","0111","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1000","0001","0000","0000","1000","0011","0000","0000","0000","0000","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0001","1010","0001","0000","0000","0000","0111","0100","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1001","0001","0000","0000","1001","0100","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1010","0001","0000","0000","0000","0111","0011","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1000","0011","0000","0001","1001","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","1001","0011","0000","0000","0001","1001","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","1001","0110","0111","1001","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0111","0111","0011","0010","0110","1000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0100","0111","0111","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","1000","1011","1011","1001","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0011","0011","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000");
signal image_G: data:=("0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0011","0100","0100","0100","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0100","1001","1100","1101","1101","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1001","1001","1001","1001","1001","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0011","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0100","1011","1010","0111","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1001","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1101","1011","0110","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1010","1010","0100","0011","0011","0011","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0110","1000","1101","0101","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0101","1100","0100","0010","0010","0001","0001","0001","0001","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","1000","1011","0100","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0111","1010","0011","0010","0010","0001","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0011","1010","0111","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1001","0111","0010","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0011","0111","1010","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0010","1001","0111","0010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0110","1011","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0010","1001","0111","0010","0010","0001","0000","0000","0000","0000","0000","0000","0001","0100","0111","1010","1010","1001","0101","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0001","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0010","0110","1011","0011","0001","0000","0000","0000","0000","0000","0000","0000","0001","0010","1001","0111","0010","0001","0000","0000","0000","0000","0000","0000","0011","0111","1011","1000","0101","0100","0110","1010","1001","0100","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0001","0110","1011","1011","0111","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","0111","1000","0111","0011","0000","0000","0000","0000","0001","0011","0101","0101","0011","0000","0000","0000","0000","0000","0000","0000","0101","1001","1001","1001","1010","1001","1010","1010","1010","1010","1000","0011","0000","0000","0000","0000","0010","0101","1011","0011","0001","0000","0000","0000","0000","0000","0000","0000","0001","0010","1001","1000","0010","0010","0000","0000","0000","0000","0000","0011","1001","0110","0010","0000","0000","0000","0000","0001","0101","1001","0101","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0110","1000","0100","0011","1000","0100","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0001","1000","0111","0101","0111","1000","0001","0000","0000","0000","0100","1001","0111","0111","1001","0011","0000","0000","0000","0000","0000","0101","1001","0100","0100","0011","0100","0100","0011","0100","0100","0011","0110","1010","0001","0000","0000","0000","0010","0101","1011","0011","0001","0000","0000","0000","0000","0000","0000","0000","0001","0010","1001","1000","0011","0010","0001","0000","0000","0000","0010","1010","0101","0001","0000","0000","0000","0000","0000","0000","0001","0100","1010","0100","0000","0000","0000","0000","0000","0000","0000","0000","0001","1001","0011","0000","0000","0011","1001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","1001","0001","0000","0010","1001","0011","0000","0000","0001","0111","0101","0000","0001","0111","0100","0000","0000","0001","0000","0000","1001","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1001","0010","0000","0000","0000","0010","0101","1011","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0010","1000","1000","0011","0010","0000","0000","0000","0001","1000","0101","0000","0000","0000","0000","0011","0010","0001","0000","0000","0000","0011","1001","0011","0000","0000","0000","0000","0000","0000","0000","0100","1000","0000","0000","0000","0001","1001","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1000","0000","0000","0000","0110","0110","0000","0000","0010","1001","0010","0000","0000","0101","0110","0001","0000","0000","0000","0000","1010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1010","0010","0000","0000","0000","0010","0101","1011","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0010","1000","1000","0011","0010","0000","0000","0000","0011","1000","0001","0000","0000","0010","1000","1010","1010","1001","0011","0000","0000","0000","0100","1001","0010","0000","0000","0000","0000","0000","0000","1000","0100","0000","0000","0000","0000","0110","0110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0101","0110","0000","0000","0000","0010","1001","0000","0000","0100","0111","0000","0000","0000","0011","1000","0001","0000","0000","0000","0001","1010","0000","0000","0000","0011","0101","0110","0110","0111","0110","0110","1000","1000","0000","0000","0000","0000","0001","0101","1011","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0010","1000","1000","0011","0001","0000","0000","0000","0111","0100","0000","0000","0001","1000","1000","0011","0011","0101","1010","0010","0000","0000","0001","1001","0011","0000","0000","0000","0000","0000","0010","1010","0010","0000","0000","0000","0000","0011","1001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0111","0101","0000","0000","0000","0001","1001","0010","0000","0111","0100","0000","0000","0000","0010","1010","0001","0000","0000","0000","0001","1010","0001","0000","0000","1000","1001","1001","1001","1001","1000","1000","1000","0001","0000","0000","0000","0000","0001","0101","1011","0100","0001","0000","0000","0000","0000","0000","0000","0000","0001","0010","1000","1000","0011","0001","0000","0000","0001","1001","0010","0000","0000","0101","0111","0001","0000","0000","0001","0110","0110","0000","0000","0000","1000","0011","0000","0000","0000","0000","0000","0110","0111","0000","0000","0000","0000","0000","0001","1001","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","1001","0010","0000","0000","0000","0000","0110","0110","0010","1001","0010","0000","0000","0000","0001","1001","0011","0000","0000","0000","0000","1011","0000","0000","0000","1010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0101","1100","0011","0001","0000","0000","0000","0000","0000","0000","0000","0001","0010","1000","1000","0011","0001","0000","0000","0001","1001","0010","0000","0000","0111","0010","0000","0000","0000","0000","0011","1001","0010","0000","0010","1010","0011","0000","0000","0000","0000","0001","1010","0011","0000","0000","0010","0010","0000","0000","0100","0111","0000","0000","0000","0000","0000","0000","0000","0000","0010","1001","0001","0000","0000","0000","0000","0011","1000","0100","1000","0000","0000","0000","0000","0000","1000","0100","0000","0000","0000","0000","1010","0001","0000","0000","1011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0101","1100","0011","0001","0000","0000","0000","0000","0000","0000","0000","0001","0010","1000","1000","0011","0010","0000","0000","0001","1010","0010","0000","0000","0111","0011","0000","0000","0000","0000","0000","0111","1000","0111","1001","0110","0000","0000","0000","0000","0000","0011","1000","0000","0000","0001","1010","1001","0001","0000","0010","1010","0010","0000","0000","0000","0000","0000","0000","0000","0011","1000","0000","0000","0000","0000","0000","0001","1000","1001","0100","0000","0000","0000","0000","0000","0100","0110","0000","0000","0000","0001","1010","0000","0000","0000","1010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0101","1100","0011","0001","0000","0000","0000","0000","0000","0000","0000","0001","0010","1000","1000","0011","0010","0000","0000","0001","1010","0001","0000","0000","0111","0010","0000","0000","0000","0001","0000","0000","0100","0101","0100","0010","0000","0000","0000","0000","0001","0111","0101","0000","0000","0011","1000","1010","0011","0000","0000","0111","0101","0000","0000","0000","0000","0000","0000","0000","0101","0110","0000","0000","0000","0000","0000","0000","0011","0110","0001","0000","0000","0000","0000","0000","0010","1000","0001","0000","0000","0001","1010","0000","0000","0000","1001","1001","1001","1000","0111","1000","0100","0000","0000","0000","0000","0000","0000","0001","0101","1100","0011","0001","0000","0000","0000","0000","0000","0000","0000","0001","0010","1000","1001","0011","0010","0000","0000","0001","1010","0001","0000","0000","0111","0010","0000","0000","0010","0011","0011","0011","0010","0010","0001","0000","0000","0000","0000","0000","0010","1010","0010","0000","0000","0111","0101","0101","0111","0000","0000","0011","1001","0000","0000","0000","0000","0000","0000","0000","0111","0100","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0001","1001","0010","0000","0000","0001","1010","0001","0000","0000","0010","0101","0110","0111","0111","1000","1011","0100","0000","0000","0000","0000","0000","0001","0101","1100","0100","0010","0000","0000","0000","0000","0000","0000","0000","0001","0010","1000","1001","0011","0001","0000","0000","0001","1010","0001","0000","0000","0111","0010","0000","0011","1001","1010","1010","1010","1010","1010","1000","0011","0000","0000","0000","0001","0101","0111","0001","0000","0001","1001","0001","0001","1001","0001","0000","0001","1010","0011","0000","0000","0000","0000","0000","0001","1001","0010","0000","0000","0010","0100","0000","0000","0000","0000","0000","0000","0001","0101","0000","0000","0001","1010","0010","0000","0000","0001","1010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","1000","0000","0000","0000","0000","0000","0001","0101","1100","0100","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","1000","1001","0011","0010","0000","0000","0001","1010","0001","0000","0000","0111","0010","0000","1000","0101","0001","0001","0001","0001","0010","0101","1001","0001","0000","0000","0001","1001","0100","0000","0000","0101","0111","0001","0001","1000","0011","0000","0000","0110","0110","0000","0000","0000","0000","0000","0010","1010","0001","0000","0001","1000","1010","0010","0000","0000","0000","0000","0001","0111","1011","0010","0000","0000","1000","0101","0000","0000","0001","1010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0100","1000","0000","0000","0000","0000","0000","0001","0100","1011","0100","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","1000","1001","0011","0010","0000","0000","0001","1010","0001","0000","0000","0111","0010","0000","1001","0011","0000","0000","0000","0000","0000","0001","1000","0011","0000","0000","0011","1001","0000","0000","0000","0101","1001","1001","1000","1010","0101","0000","0000","0010","1001","0001","0000","0000","0000","0000","0011","1001","0001","0000","0001","1010","0110","0101","0000","0000","0000","0000","0001","1010","0111","0100","0000","0000","0110","0111","0000","0000","0001","1010","0000","0000","0000","0001","0011","0011","0011","0010","0011","1001","0101","0000","0000","0000","0000","0000","0001","0100","1011","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0010","1000","1001","0011","0001","0001","0000","0010","1010","0001","0000","0000","0111","0010","0000","0111","1000","0100","0011","0001","0000","0000","0000","0111","0011","0000","0000","0111","0101","0000","0000","0000","0001","0100","0101","0101","0101","0010","0000","0000","0000","1000","0011","0000","0000","0000","0000","0101","0111","0000","0000","0011","1001","0011","1000","0001","0000","0000","0000","0011","1000","0101","0111","0000","0000","0010","1001","0000","0000","0001","1010","0000","0000","0000","1000","1001","1001","1010","1010","1001","1001","0000","0000","0000","0000","0000","0000","0001","0100","1100","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0010","1000","1001","0011","0010","0000","0000","0001","1010","0001","0000","0000","1000","0001","0000","0010","1000","1010","1010","1000","0000","0000","0000","1000","0011","0000","0001","1001","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0101","0111","0000","0000","0000","0000","0110","0100","0000","0000","0101","0111","0001","1001","0010","0000","0000","0000","0111","0101","0010","1001","0000","0000","0001","1001","0001","0000","0001","1001","0000","0000","0000","1011","0010","0000","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0001","0100","1100","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0010","1000","1001","0011","0001","0000","0000","0001","1010","0010","0000","0000","0110","0101","0000","0000","0000","0001","0011","1000","0001","0000","0001","1001","0010","0000","0100","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","1010","0001","0000","0000","0000","1000","0010","0000","0000","0110","0100","0000","0111","0100","0000","0000","0001","1001","0010","0001","1010","0001","0000","0000","1000","0010","0000","0001","1010","0000","0000","0001","1010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0100","1100","0100","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","1000","1001","0010","0001","0000","0000","0000","1000","0100","0000","0000","0010","1010","0110","0001","0001","0010","1001","0100","0000","0000","0001","1001","0001","0000","0111","0100","0000","0000","0010","1000","1000","0111","0111","1000","0111","0111","0101","0000","0000","0000","0111","0100","0000","0000","0001","1001","0001","0000","0000","1000","0011","0000","0011","1001","0110","0100","1000","0111","0000","0000","1001","0010","0000","0000","0111","0011","0000","0001","1010","0000","0000","0001","1011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0100","1100","0100","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","0111","1001","0011","0010","0000","0000","0000","0101","1000","0001","0000","0000","0010","1001","1011","1010","1011","0110","0000","0000","0000","0101","0111","0000","0001","1001","0001","0000","0000","0110","1000","0110","0110","0110","0110","0111","1000","1010","0011","0000","0000","0011","1000","0001","0000","0010","1001","0001","0000","0000","1001","0001","0000","0000","0100","1010","1011","1000","0001","0000","0000","0111","0011","0000","0000","0101","0101","0000","0001","1001","0000","0000","0000","1001","0011","0010","0010","0010","0010","0001","0010","0000","0000","0000","0000","0000","0001","0100","1100","0100","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","0111","1001","0011","0010","0000","0000","0000","0001","1001","0101","0000","0000","0000","0010","0100","0100","0011","0000","0000","0000","0011","1001","0010","0000","0101","0111","0000","0000","0010","1001","0011","0000","0000","0001","0000","0000","0001","0101","0110","0000","0000","0001","1010","0010","0000","0101","1000","0000","0000","0001","1001","0001","0000","0000","0000","0001","0001","0001","0000","0000","0000","0110","0011","0000","0000","0011","1000","0000","0000","1010","0000","0000","0000","0101","1010","1010","1010","1001","1010","1010","1001","0101","0000","0000","0000","0000","0001","0100","1100","0100","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","0111","1001","0011","0010","0000","0000","0000","0000","0011","1010","0011","0000","0000","0000","0000","0000","0000","0000","0000","0001","1000","0110","0000","0000","1000","0100","0000","0000","0011","1000","0000","0000","0000","0000","0000","0000","0000","0010","1010","0010","0000","0000","0111","0100","0000","0110","0101","0000","0000","0100","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0101","0101","0000","0000","0010","1010","0001","0000","1001","0000","0000","0000","0000","0001","0001","0001","0010","0010","0001","0011","1010","0001","0000","0000","0000","0001","0100","1100","0100","0010","0000","0000","0000","0000","0000","0000","0000","0001","0010","0111","1001","0011","0010","0000","0000","0000","0000","0001","0100","1010","0100","0010","0000","0000","0000","0000","0001","0011","1001","1000","0001","0000","0000","0111","0101","0000","0001","0111","0110","0000","0000","0000","0000","0000","0000","0000","0001","1000","0101","0000","0001","1000","0100","0000","0110","0101","0000","0001","0110","0110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1000","0001","0000","0001","1010","0001","0000","1010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1001","0001","0000","0000","0000","0001","0100","1100","0100","0010","0000","0000","0000","0000","0000","0000","0000","0000","0010","0111","1001","0011","0010","0000","0000","0000","0000","0000","0000","0011","1001","1001","0111","0111","0110","0110","1000","1001","0110","0001","0000","0000","0000","0011","1001","0111","1000","0111","0010","0000","0000","0000","0000","0000","0000","0000","0000","0100","1001","0110","0110","1001","0010","0000","0010","1010","0111","0111","1001","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1001","0110","0011","0111","1001","0001","0000","1001","0110","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","1010","0000","0000","0000","0000","0001","0100","1100","0100","0010","0001","0000","0000","0000","0000","0000","0000","0000","0010","0111","1001","0011","0010","0000","0000","0000","0000","0000","0000","0000","0010","0100","0110","0111","1000","0111","0100","0010","0000","0000","0000","0000","0000","0001","0011","0111","0100","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0100","0111","1000","0011","0000","0000","0000","0011","0111","0110","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1001","1011","1001","0011","0000","0000","0010","1011","1011","1100","1011","1100","1011","1011","1011","1011","1011","1100","0111","0000","0000","0000","0000","0001","0100","1100","0100","0010","0001","0000","0000","0000","0000","0000","0000","0000","0010","0111","1001","0011","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0000","0000","0000","0000","0001","0011","0011","0100","0100","0100","0100","0100","0101","0101","0100","0000","0000","0000","0000","0000","0001","0100","1100","0100","0010","0001","0000","0000","0000","0000","0000","0000","0000","0010","0111","1001","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0100","1100","0100","0010","0001","0000","0000","0000","0000","0000","0000","0000","0010","0111","1010","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0011","0011","0010","0001","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0100","1101","0100","0010","0001","0000","0000","0000","0000","0000","0000","0000","0001","0111","1010","0011","0001","0000","0000","0000","0000","0000","0000","0000","0011","1000","1001","1001","1010","1010","1001","1001","1000","0011","0000","0000","0000","0000","0000","0001","0111","1001","0111","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0111","1000","0100","0000","0000","0000","0001","0100","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0011","0000","0000","0000","0001","0101","0111","0111","0111","0111","0111","0111","0110","0101","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0100","1101","0100","0010","0001","0000","0000","0000","0000","0000","0000","0000","0001","0111","1010","0011","0001","0000","0000","0000","0000","0000","0000","0101","1010","0110","0010","0001","0001","0001","0001","0011","0110","1011","0101","0000","0000","0000","0000","0110","1000","0100","1000","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1010","0111","0110","1011","0010","0000","0000","0100","1010","0101","0100","0100","0100","0100","0100","0101","0101","0100","0101","0111","1001","0001","0000","0000","0110","1001","0101","0101","0100","0101","0110","0101","0110","0111","1010","1000","0011","0001","0000","0000","0000","0000","0000","0000","0001","0100","1100","0100","0010","0001","0000","0000","0000","0000","0000","0000","0000","0001","0111","1010","0011","0010","0000","0000","0000","0000","0000","0100","1011","0011","0000","0000","0000","0000","0000","0000","0000","0000","0011","1011","0101","0000","0000","0000","1001","0001","0000","0000","1010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","1001","0000","0000","0100","1000","0000","0010","1001","0100","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1000","0011","0000","0000","1000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0001","0111","1010","0101","0000","0000","0000","0000","0000","0000","0001","0011","1100","0100","0010","0001","0000","0000","0000","0000","0000","0000","0000","0010","0111","1010","0011","0001","0000","0000","0000","0000","0100","1010","0011","0000","0000","0000","0000","0001","0001","0000","0000","0000","0000","0010","1010","0100","0000","0000","1001","0001","0000","0000","0111","0110","0000","0000","0000","0000","0000","0000","0000","0000","0000","1000","0011","0000","0000","0011","0111","0000","0010","1001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1001","0011","0000","0001","1001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","1010","0100","0000","0000","0000","0000","0000","0001","0011","1100","0100","0010","0001","0000","0000","0000","0000","0000","0000","0000","0010","0111","1010","0011","0001","0000","0000","0000","0000","1001","0100","0000","0000","0000","0010","1001","1100","1100","1001","0100","0000","0000","0000","0100","1010","0000","0000","1000","0011","0000","0000","0011","1010","0000","0000","0000","0000","0000","0000","0000","0000","0001","1010","0000","0000","0000","0111","0100","0000","0010","1000","0000","0000","0000","0010","0011","0010","0010","0010","0010","0010","0010","0011","1010","0001","0000","0000","1010","0010","0000","0000","0011","0100","0100","0011","0010","0001","0000","0000","0000","0100","1001","0001","0000","0000","0000","0000","0001","0011","1100","0100","0010","0001","0000","0000","0000","0000","0000","0000","0000","0010","0111","1010","0010","0001","0000","0000","0000","0100","1001","0000","0000","0000","0101","1010","0111","0100","0100","0110","1010","0110","0000","0000","0000","0111","0101","0000","0101","1000","0000","0000","0001","1001","0001","0000","0000","0000","0000","0000","0000","0000","0101","1000","0000","0000","0001","1010","0000","0000","0010","1000","0000","0000","0001","0111","1010","1011","1011","1010","1011","1010","1011","1010","0100","0001","0000","0001","1001","0001","0000","0001","1001","1001","1010","1010","1010","1000","0011","0000","0000","0000","1001","0011","0000","0000","0000","0000","0001","0011","1100","0100","0010","0001","0000","0000","0000","0000","0000","0000","0000","0010","0111","1010","0011","0001","0000","0000","0000","1001","0011","0000","0000","0011","1010","0011","0000","0000","0000","0000","0010","1001","0100","0000","0000","0010","1001","0000","0001","1010","0001","0000","0000","0110","0101","0000","0000","0000","0000","0000","0000","0000","1001","0011","0000","0000","0101","1000","0000","0000","0011","1000","0000","0000","0010","1010","0011","0001","0010","0010","0010","0010","0010","0010","0000","0000","0000","0001","1010","0001","0000","0001","1001","0010","0000","0001","0010","0101","1010","0001","0000","0000","0100","1000","0000","0000","0000","0000","0001","0011","1100","0100","0010","0001","0000","0000","0000","0000","0000","0000","0000","0010","0110","1010","0010","0001","0000","0000","0000","1010","0001","0000","0000","1001","0100","0000","0000","0000","0000","0000","0000","0100","1001","0000","0000","0001","1001","0001","0000","1000","0100","0000","0000","0011","1010","0000","0000","0000","0000","0000","0000","0010","1010","0000","0000","0000","1001","0100","0000","0000","0011","1000","0000","0000","0001","1010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1001","0001","0000","0000","1001","0001","0000","0000","0000","0001","0111","0011","0000","0000","0010","1010","0001","0000","0000","0000","0001","0011","1100","0101","0010","0001","0000","0000","0000","0000","0000","0000","0000","0010","0110","1010","0010","0001","0000","0000","0001","1010","0001","0000","0000","1001","0001","0000","0000","0000","0000","0000","0000","0001","1001","0000","0000","0000","1010","0001","0000","0100","1000","0000","0000","0000","1010","0011","0000","0000","0000","0000","0000","0110","0111","0000","0000","0010","1011","0000","0000","0000","0011","1000","0000","0000","0001","1010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1010","0001","0000","0001","1001","0010","0000","0000","0000","0000","0110","0101","0000","0000","0001","1001","0001","0000","0000","0000","0001","0011","1100","0101","0010","0001","0000","0000","0000","0000","0000","0000","0001","0010","0110","1010","0010","0001","0000","0000","0001","1011","0000","0000","0000","1010","0000","0000","0000","0000","0000","0000","0000","0010","1010","0000","0000","0000","1010","0000","0000","0000","1010","0010","0000","0000","0110","0110","0000","0000","0000","0000","0001","1010","0010","0000","0000","0110","0111","0000","0000","0000","0011","1000","0000","0000","0010","1001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1001","0010","0000","0000","1000","0001","0000","0000","0000","0000","0101","0101","0000","0000","0001","1001","0001","0000","0000","0000","0001","0011","1100","0101","0010","0001","0000","0000","0000","0000","0000","0000","0001","0010","0110","1010","0011","0001","0000","0000","0001","1011","0000","0000","0000","1010","0000","0000","0000","0000","0000","0000","0000","0001","1010","0000","0000","0001","1010","0001","0000","0000","1000","0101","0000","0000","0011","1001","0000","0000","0000","0000","0100","1001","0000","0000","0000","1010","0010","0000","0000","0000","0011","1000","0000","0000","0001","1010","0010","0010","0010","0010","0010","0001","0000","0000","0000","0000","0000","0001","1010","0001","0000","0001","1001","0001","0000","0000","0000","0010","1001","0011","0000","0000","0010","1010","0001","0000","0000","0000","0001","0011","1100","0101","0010","0001","0000","0000","0000","0000","0000","0000","0000","0010","0110","1010","0010","0001","0000","0000","0001","1011","0000","0000","0000","1010","0000","0000","0000","0000","0000","0000","0000","0001","1010","0000","0000","0000","1010","0001","0000","0000","0011","1001","0000","0000","0000","1001","0010","0000","0000","0000","0111","0101","0000","0000","0011","1001","0000","0000","0000","0000","0011","1000","0000","0000","0001","0111","1001","1001","1001","1001","1001","1001","1000","0001","0000","0000","0000","0001","1010","0001","0000","0001","1001","0100","0010","0011","0100","1001","1000","0001","0000","0000","0011","1001","0000","0000","0000","0000","0000","0011","1100","0101","0010","0001","0000","0000","0000","0000","0000","0000","0000","0010","0110","1011","0010","0001","0000","0000","0001","1011","0000","0000","0001","1011","0000","0000","0000","0000","0000","0000","0000","0001","1010","0000","0000","0000","1010","0001","0000","0000","0001","1011","0001","0000","0000","0110","0110","0000","0000","0000","1011","0010","0000","0000","0111","0101","0000","0000","0000","0000","0011","1000","0000","0000","0000","0001","0010","0010","0010","0010","0011","0011","1001","0100","0000","0000","0000","0001","1010","0001","0000","0001","1001","1011","1100","1100","1011","0111","0010","0000","0000","0000","0110","0110","0000","0000","0000","0000","0000","0011","1100","0101","0010","0001","0000","0000","0000","0000","0000","0000","0000","0010","0110","1011","0011","0001","0000","0000","0001","1011","0000","0000","0001","1011","0001","0000","0000","0000","0000","0000","0000","0001","1010","0000","0000","0000","1010","0001","0000","0000","0000","0111","0110","0000","0000","0010","1010","0000","0000","0100","1000","0000","0000","0001","1010","0010","0000","0000","0000","0000","0011","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0101","0111","0000","0000","0000","0001","1001","0001","0000","0000","0010","0010","0010","0010","0010","0001","0000","0000","0000","0010","1010","0010","0000","0000","0000","0000","0000","0011","1100","0101","0010","0001","0000","0000","0000","0000","0000","0000","0000","0010","0110","1011","0011","0001","0000","0000","0001","1011","0000","0000","0001","1011","0001","0000","0000","0000","0000","0000","0000","0001","1010","0000","0000","0000","1010","0001","0000","0000","0000","0010","1001","0000","0000","0000","1010","0011","0000","1000","0011","0000","0000","0100","1001","0000","0000","0000","0000","0000","0011","1000","0001","0000","0001","0000","0000","0000","0000","0000","0000","0000","0110","0110","0000","0000","0000","0001","1001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0111","0110","0000","0000","0000","0000","0000","0001","0011","1100","0101","0010","0001","0000","0000","0000","0000","0000","0000","0000","0010","0110","1011","0011","0001","0000","0000","0001","1011","0000","0000","0001","1011","0001","0000","0000","0000","0000","0000","0000","0001","1001","0000","0000","0000","1011","0001","0000","0000","0000","0000","1010","0010","0000","0000","0101","0111","0001","1010","0001","0000","0000","1000","0100","0000","0000","0000","0000","0000","0011","1000","0000","0000","0001","0011","0100","0100","0100","0100","0100","0101","1001","0010","0000","0000","0000","0001","1010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","1011","0010","0000","0000","0000","0000","0000","0001","0011","1100","0101","0010","0001","0000","0000","0000","0000","0000","0000","0000","0010","0110","1011","0011","0001","0000","0000","0001","1011","0000","0000","0000","1011","0001","0000","0000","0000","0000","0000","0000","0001","1001","0000","0000","0000","1011","0001","0000","0000","0000","0000","0110","0110","0000","0000","0001","1010","0111","1000","0000","0000","0001","1010","0001","0000","0000","0000","0000","0000","0011","1000","0000","0000","0001","1001","0111","0111","0111","1000","1000","0111","0101","0000","0000","0000","0000","0001","1010","0001","0000","0000","0011","0101","0101","0101","0110","0101","0000","0000","0001","0111","0110","0000","0000","0000","0000","0000","0001","0011","1100","0101","0010","0001","0000","0000","0000","0000","0000","0000","0000","0010","0110","1011","0011","0001","0000","0000","0001","1011","0000","0000","0001","1010","0000","0000","0000","0000","0000","0000","0000","0001","1001","0000","0000","0000","1011","0001","0000","0000","0000","0000","0001","1010","0000","0000","0000","0110","1010","0010","0000","0000","0101","1000","0000","0000","0000","0000","0000","0000","0011","1000","0000","0000","0001","1010","0001","0000","0000","0001","0001","0001","0000","0000","0000","0000","0000","0001","1010","0001","0000","0000","1000","1000","1000","1000","1000","1010","0011","0000","0000","0010","1001","0010","0000","0000","0000","0000","0001","0011","1100","0110","0010","0001","0000","0000","0000","0000","0000","0000","0000","0010","0110","1011","0011","0001","0000","0000","0001","1011","0000","0000","0001","1010","0000","0000","0000","0000","0000","0000","0000","0010","1001","0000","0000","0000","1011","0001","0000","0000","0000","0000","0000","1001","0010","0000","0000","0001","0010","0000","0000","0000","1001","0011","0000","0000","0000","0000","0000","0000","0011","1000","0000","0000","0001","1010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1010","0001","0000","0001","1001","0001","0000","0001","0000","0101","1000","0001","0000","0001","1001","0010","0000","0000","0000","0000","0001","0011","1100","0110","0010","0001","0000","0000","0000","0000","0000","0000","0000","0010","0110","1011","0011","0001","0000","0000","0000","1011","0000","0000","0000","1000","0100","0000","0000","0000","0000","0000","0000","1000","0101","0000","0000","0001","1010","0000","0000","0000","0000","0000","0000","0110","0111","0000","0000","0000","0000","0000","0000","0001","1010","0000","0000","0000","0000","0000","0000","0000","0011","1000","0000","0000","0010","1010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1010","0001","0000","0001","1001","0001","0000","0000","0000","0001","1010","0001","0000","0000","1000","0010","0000","0000","0000","0000","0000","0011","1100","0110","0010","0001","0000","0000","0000","0000","0000","0000","0000","0010","0110","1011","0011","0001","0000","0000","0000","1010","0010","0000","0000","0011","1010","0011","0000","0000","0000","0000","0110","1010","0001","0000","0000","0011","1001","0000","0000","0000","0000","0000","0000","0010","1010","0001","0000","0000","0000","0000","0000","0110","0110","0000","0000","0000","0000","0000","0000","0000","0011","1000","0000","0000","0001","1010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1010","0001","0000","0001","1001","0001","0000","0000","0000","0001","1001","0010","0000","0000","1000","0010","0000","0000","0000","0000","0000","0011","1100","0110","0010","0001","0000","0000","0000","0000","0000","0000","0000","0010","0110","1011","0011","0001","0000","0000","0000","0110","0111","0000","0000","0000","0101","1010","0110","0100","0101","1000","1001","0010","0000","0000","0000","1000","0101","0000","0000","0000","0000","0000","0000","0000","1001","0011","0000","0000","0000","0000","0000","1010","0010","0000","0000","0000","0000","0000","0000","0000","0010","1000","0000","0000","0010","1010","0011","0010","0010","0010","0001","0010","0001","0010","0000","0000","0000","0001","1010","0001","0000","0001","1000","0001","0000","0000","0000","0001","1001","0010","0000","0000","1000","0011","0000","0000","0000","0000","0001","0011","1100","0110","0010","0001","0000","0000","0000","0000","0000","0000","0000","0001","0101","1011","0011","0001","0000","0000","0000","0001","1011","0011","0000","0000","0000","0100","0111","1001","1000","0110","0001","0000","0000","0000","0101","1001","0001","0000","0000","0000","0000","0000","0000","0000","0101","0111","0000","0000","0000","0000","0011","1001","0000","0000","0000","0000","0000","0000","0000","0000","0011","1000","0000","0000","0001","1000","1011","1011","1011","1010","1011","1010","1010","1001","0011","0000","0000","0010","1010","0001","0000","0000","1001","0001","0000","0000","0000","0001","1001","0010","0000","0000","0111","0100","0000","0000","0000","0000","0001","0011","1011","0110","0010","0001","0000","0000","0000","0000","0000","0000","0000","0001","0101","1011","0011","0001","0000","0001","0000","0000","0101","1011","0011","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0011","1010","0011","0000","0000","0000","0000","0000","0000","0000","0000","0010","1011","0000","0000","0000","0000","1000","0110","0000","0000","0000","0000","0000","0000","0000","0000","0011","0111","0000","0000","0000","0010","0011","0011","0011","0100","0100","0101","0100","0110","1010","0001","0000","0001","1001","0001","0000","0001","1000","0001","0000","0000","0000","0001","1001","0010","0000","0000","0110","0100","0000","0000","0000","0000","0001","0011","1011","0110","0010","0001","0000","0000","0000","0000","0000","0000","0000","0001","0101","1100","0011","0010","0000","0000","0000","0000","0000","0100","1010","0100","0000","0000","0000","0000","0000","0000","0000","0001","0101","1001","0100","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1001","0100","0000","0000","0001","1010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0011","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1001","0010","0000","0001","1010","0001","0000","0000","1001","0010","0000","0000","0000","0001","1001","0001","0000","0000","0111","0101","0000","0000","0000","0000","0000","0011","1011","0110","0010","0001","0000","0000","0000","0000","0000","0000","0000","0001","0101","1100","0011","0010","0000","0000","0000","0000","0000","0000","0100","1011","0111","0010","0001","0000","0000","0000","0011","1000","1011","0100","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","1001","0010","0001","0110","1000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0010","1010","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0001","1010","0010","0000","0001","1001","0001","0000","0001","1001","0001","0000","0000","0000","0000","1000","0010","0000","0000","0111","0100","0000","0000","0000","0000","0000","0011","1011","0110","0010","0001","0000","0000","0000","0000","0000","0000","0000","0001","0101","1100","0011","0001","0001","0000","0000","0000","0000","0000","0000","0010","1001","1010","1001","1001","1001","1001","1010","1000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1000","1010","1010","1010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0111","1001","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","1000","1000","0001","0000","0000","1000","0111","0101","1000","0111","0000","0000","0000","0000","0000","0101","1000","0100","0110","1010","0010","0000","0000","0000","0000","0000","0011","1011","0110","0010","0001","0000","0000","0000","0000","0000","0000","0000","0001","0101","1100","0011","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0011","0100","0100","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0010","0000","0000","0000","0010","0101","0110","0101","0001","0000","0000","0000","0000","0000","0001","0101","0111","0110","0011","0000","0000","0000","0000","0000","0000","0011","1011","0111","0010","0001","0000","0000","0000","0000","0000","0000","0000","0001","0100","1100","0100","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0001","0000","0000","0000","0000","0000","0000","0000","0011","1011","0110","0011","0001","0000","0000","0000","0000","0000","0000","0000","0001","0011","1011","0111","0010","0010","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0011","1100","0101","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0010","0111","1100","0110","0011","0011","0011","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0010","0001","0010","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0001","0001","0001","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0001","0001","0001","0000","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0010","0101","1101","0100","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0011","1001","1100","1001","0110","0101","0100","0010","0001","0000","0001","0011","0011","0011","0000","0000","0000","0001","0011","0100","0011","0011","0011","0011","0011","0100","0011","0011","0100","0010","0000","0000","0000","0001","0010","0011","0011","0010","0001","0000","0000","0001","0010","0011","0010","0010","0010","0010","0010","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0000","0000","0000","0001","0010","0001","0001","0000","0000","0000","0000","0001","0001","0001","0010","0100","1001","1010","0100","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0011","0111","1001","1011","1100","1011","0110","0001","0001","0011","0111","1011","1000","0011","0000","0000","0011","1001","1011","1011","1100","1100","1011","1100","1011","1100","1100","1011","0111","0001","0000","0001","0010","0111","1010","1001","0101","0001","0001","0000","0010","0110","1000","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0110","0011","0001","0000","0010","0100","0110","0101","0001","0001","0000","0000","0000","0010","0101","0110","0110","1010","1011","0101","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0010","0011","0101","0110","1001","1001","0010","0001","0100","1110","1001","1101","0110","0001","0010","0101","1100","1001","1000","1000","1000","1000","1000","1000","1000","1000","1001","1100","0100","0001","0001","0110","1101","1010","1011","1100","0100","0000","0010","0110","1101","1100","1011","1011","1011","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1101","1101","1100","1101","1101","1101","1101","1101","1101","1110","0110","0001","0001","0100","1101","1110","1101","0110","0010","0000","0000","0001","0101","1101","1110","1110","1010","0101","0011","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0010","0011","0110","1011","0010","0010","0110","1010","0100","1000","1001","0010","0010","0110","1011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","1011","0100","0001","0011","1010","1000","0100","0101","1011","0110","0010","0001","1000","1000","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0111","1010","0010","0010","0111","1010","0101","1001","1010","0010","0001","0000","0001","1000","1001","0101","0100","0100","0010","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0101","1011","0011","0010","0110","1010","0011","0111","1010","0011","0011","0110","1011","0011","0010","0001","0001","0001","0001","0010","0001","0010","0011","1011","0100","0010","0011","1011","0111","0010","0011","1010","0111","0010","0010","1000","1000","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0101","1011","0011","0010","1000","1001","0011","0101","1100","0011","0001","0000","0010","1001","0111","0011","0010","0010","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0110","1010","0011","0010","0111","1010","0011","0101","1100","0100","0100","1000","1010","0010","0001","0001","0000","0001","0001","0001","0001","0010","0011","1011","0100","0010","0011","1011","0110","0011","0011","1010","0111","0010","0010","1000","1000","0011","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0101","1100","0011","0011","1001","1000","0011","0101","1100","0011","0001","0000","0010","1001","0111","0011","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0101","1011","0011","0011","0111","1010","0011","0100","1011","1011","1011","1100","0111","0001","0000","0000","0000","0000","0000","0000","0001","0001","0011","1011","0101","0010","0011","1011","0110","0010","0011","1001","1000","0010","0011","1000","1000","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0010","0100","1100","0100","0100","1010","1000","0010","0101","1100","0011","0001","0000","0010","1001","0111","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0101","1011","0011","0010","0111","1010","0011","0010","0100","0111","1000","0110","0011","0001","0000","0000","0000","0000","0000","0000","0000","0001","0011","1011","0101","0010","0011","1011","0110","0010","0011","1001","1000","0011","0011","1001","1000","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0011","1011","1011","1010","1101","0101","0010","0100","1100","0011","0001","0001","0010","1001","0110","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0110","1010","0100","0011","0111","1010","0011","0001","0010","0010","0011","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0011","1011","0101","0010","0011","1011","0110","0010","0010","1000","1001","0100","0100","1010","0111","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0101","1010","1011","0110","0010","0010","0100","1100","0011","0001","0001","0011","1001","0110","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0110","1011","0011","0011","1000","1001","0010","0000","0001","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0011","1011","0101","0010","0011","1011","0110","0010","0010","0101","1100","1010","1010","1100","0101","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0010","0011","0011","0010","0010","0010","0100","1100","0011","0001","0001","0011","1001","0110","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0101","1100","0111","0110","1011","0111","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0011","1011","0101","0010","0011","1011","0110","0001","0001","0011","0110","1010","1011","0110","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0010","0010","0001","0001","0010","0100","1100","0100","0010","0001","0011","1001","0110","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","1000","1100","1100","1010","0100","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0011","1011","0101","0011","0011","1011","0110","0010","0001","0001","0010","0011","0011","0010","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0000","0001","0100","1101","0100","0010","0001","0011","1001","0110","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0100","0100","0011","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","1011","0101","0011","0011","1011","0110","0001","0000","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0100","1101","0100","0010","0010","0011","1010","0110","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0010","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","1010","0111","0100","0100","1100","0101","0001","0000","0001","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0100","1100","0101","0011","0010","0100","1100","0101","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0010","0110","1101","1010","1011","1011","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1010","1010","0110","0101","1001","1011","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","0110","1010","1001","0101","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0100","1011","1110","1110","1100","0101","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0011","0011","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0011","0101","0110","0100","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0010","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000");
signal image_B: data:=("0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0010","0010","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0011","0100","0101","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0010","0010","0011","0010","0010","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0011","0101","0111","1000","1001","1001","1001","1001","1000","1001","1001","1001","1001","1001","1001","1001","1001","1000","1001","1001","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0101","0100","0011","0001","0001","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0001","0010","0100","1000","1101","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1101","1101","1101","1101","1101","1101","1101","1101","1101","1100","1100","1100","1100","1100","1100","1100","1100","1100","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1011","1010","1010","1001","0111","0101","0011","0010","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0001","0010","0111","1111","1111","1100","1010","1010","1010","1010","1010","1010","1011","1011","1011","1011","1011","1011","1011","1011","1100","1100","1100","1100","1100","1100","1100","1100","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1110","1110","1110","1110","1110","1110","1110","1110","1110","1110","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1010","0110","0011","0001","0000","0000","0000","0000","0000","0000","0000","0001","0001","0010","0101","1101","1110","1001","0111","0110","0110","0101","0101","0110","0101","0101","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1001","1000","1000","1000","1001","1001","1001","1001","1001","1001","1001","1010","1101","1111","1001","0101","0010","0001","0000","0000","0000","0000","0000","0000","0001","0001","0010","1000","1111","1000","0111","0110","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0100","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0110","0110","0110","0110","0110","0101","0110","0110","1000","1101","1111","0111","0100","0001","0000","0000","0000","0000","0000","0000","0001","0001","0100","1010","1110","1000","0110","0101","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0010","0011","0011","0100","0100","0011","0011","0011","0100","0101","0110","1000","1111","1011","0101","0010","0001","0000","0000","0000","0000","0000","0000","0001","0100","1100","1100","0111","0101","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0000","0001","0000","0000","0000","0000","0001","0001","0010","0001","0001","0001","0001","0001","0011","0101","0111","1011","1110","0110","0011","0001","0000","0000","0000","0000","0000","0000","0001","0100","1101","1100","0111","0100","0010","0001","0000","0000","0000","0000","0000","0000","0000","0001","0010","0010","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0011","0101","1010","1111","0111","0100","0001","0000","0000","0000","0000","0000","0000","0001","0101","1101","1100","0110","0100","0010","0001","0000","0000","0000","0000","0000","0010","0100","1000","1010","1011","1010","0110","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0010","0001","0000","0000","0000","0000","0000","0000","0001","0010","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0010","0001","0001","0001","0001","0001","0010","0001","0001","0000","0000","0000","0000","0001","0010","0101","1001","1111","0111","0100","0001","0000","0000","0000","0000","0000","0000","0001","0101","1101","1100","0110","0100","0010","0001","0000","0000","0000","0001","0100","1000","1100","1001","0110","0101","0110","1011","1010","0101","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0111","1011","1100","1000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","0111","1001","0111","0100","0001","0000","0000","0000","0010","0100","0110","0110","0100","0000","0000","0000","0000","0000","0000","0000","0110","1010","1010","1010","1010","1010","1011","1010","1010","1011","1001","0011","0000","0000","0001","0010","0100","1001","1111","0111","0100","0001","0000","0000","0000","0000","0000","0000","0010","0101","1101","1100","0110","0100","0010","0001","0000","0000","0001","0101","1010","0111","0011","0001","0000","0000","0000","0001","0110","1010","0110","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0111","1001","0100","0011","1001","0110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1001","0111","0110","1000","1001","0010","0000","0000","0000","0100","1010","1000","1001","1010","0011","0000","0000","0000","0000","0000","0110","1010","0101","0101","0100","0101","0101","0100","0100","0100","0100","0110","1010","0001","0000","0000","0010","0100","1001","1111","0111","0100","0001","0000","0000","0000","0000","0000","0000","0010","0101","1101","1100","0110","0100","0010","0000","0000","0000","0011","1100","0110","0010","0000","0000","0000","0000","0000","0000","0001","0100","1011","0101","0001","0000","0000","0000","0000","0000","0000","0000","0010","1010","0011","0000","0000","0100","1010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1010","0010","0000","0010","1010","0100","0000","0000","0001","1000","0101","0000","0010","1000","0101","0000","0000","0000","0000","0001","1010","0100","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1010","0010","0000","0000","0001","0100","1001","1111","0111","0100","0001","0000","0000","0000","0000","0000","0000","0010","0101","1101","1100","0110","0100","0001","0000","0000","0010","1001","0110","0001","0000","0000","0000","0011","0010","0001","0000","0000","0000","0100","1011","0100","0000","0000","0000","0000","0000","0000","0000","0101","1001","0001","0000","0000","0010","1010","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","1001","0000","0000","0000","0111","0111","0000","0000","0010","1010","0010","0000","0000","0101","0110","0001","0000","0000","0000","0001","1011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1010","0010","0000","0000","0001","0100","1001","1111","0111","0100","0001","0000","0000","0000","0000","0000","0000","0010","0101","1101","1100","0110","0100","0001","0000","0000","0100","1010","0010","0000","0000","0011","1001","1011","1011","1010","0100","0000","0000","0000","0101","1010","0010","0000","0000","0000","0000","0000","0000","1000","0100","0000","0000","0000","0001","0110","0110","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0110","0111","0000","0000","0000","0011","1010","0000","0000","0100","1000","0000","0000","0000","0011","1001","0001","0000","0000","0000","0001","1011","0000","0000","0000","0011","0110","0111","0111","1000","0111","0111","1001","1001","0000","0000","0000","0001","0100","1001","1111","0111","0100","0001","0000","0000","0000","0000","0000","0000","0010","0110","1101","1101","0110","0011","0010","0000","0001","1000","0101","0000","0000","0010","1001","1000","0011","0011","0110","1011","0010","0000","0000","0001","1010","0011","0000","0000","0000","0000","0000","0010","1010","0010","0000","0000","0000","0000","0011","1010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0001","1000","0101","0000","0000","0000","0010","1010","0011","0000","1000","0100","0000","0000","0000","0011","1010","0010","0000","0000","0000","0001","1011","0001","0000","0001","1001","1010","1010","1010","1010","1001","1001","1001","0010","0000","0000","0000","0001","0100","1001","1111","0111","0100","0001","0000","0000","0000","0000","0000","0001","0010","0101","1101","1101","0110","0011","0001","0000","0001","1010","0011","0000","0000","0110","1001","0001","0000","0000","0001","0111","0111","0001","0000","0000","1001","0100","0000","0000","0000","0000","0001","0110","0111","0000","0000","0000","0000","0000","0001","1001","0100","0000","0000","0000","0000","0000","0000","0000","0000","0010","1011","0011","0000","0000","0000","0001","0111","0110","0010","1010","0010","0000","0000","0000","0001","1010","0100","0000","0000","0000","0001","1011","0001","0000","0001","1010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0100","1000","1111","0111","0101","0001","0000","0000","0000","0000","0000","0001","0010","0101","1101","1101","0110","0011","0001","0000","0001","1010","0011","0000","0000","1000","0011","0000","0000","0000","0000","0011","1010","0010","0001","0011","1011","0011","0000","0000","0000","0000","0010","1011","0011","0000","0000","0010","0011","0000","0000","0101","1000","0001","0000","0000","0000","0000","0000","0000","0000","0011","1011","0010","0000","0000","0000","0000","0011","1001","0101","1001","0000","0000","0000","0000","0001","1001","0101","0000","0000","0000","0001","1010","0001","0000","0000","1011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0100","1000","1111","0111","0101","0001","0000","0000","0000","0000","0000","0001","0010","0110","1101","1101","0110","0011","0001","0000","0001","1010","0010","0000","0000","1000","0100","0000","0000","0000","0000","0000","1000","1001","1000","1010","0111","0001","0000","0000","0000","0000","0100","1001","0001","0000","0010","1010","1001","0001","0000","0010","1011","0011","0000","0000","0000","0000","0000","0000","0000","0101","1001","0001","0000","0000","0000","0000","0001","1001","1010","0100","0000","0000","0000","0000","0000","0110","1000","0001","0000","0000","0001","1010","0001","0000","0000","1011","0010","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0001","0100","1000","1111","1000","0101","0001","0000","0000","0000","0000","0000","0000","0010","0110","1101","1101","0110","0011","0001","0000","0010","1011","0010","0000","0001","1000","0011","0000","0000","0000","0001","0001","0010","0101","0111","0100","0010","0000","0000","0000","0000","0001","1000","0110","0000","0000","0011","1001","1010","0011","0000","0001","1000","0110","0000","0000","0000","0000","0000","0000","0000","0110","0111","0000","0000","0000","0000","0000","0000","0100","0110","0001","0000","0000","0000","0000","0000","0011","1001","0010","0000","0000","0001","1010","0001","0000","0000","1001","1010","1001","1001","1000","1001","0101","0001","0000","0000","0000","0000","0001","0100","1000","1111","1000","0101","0001","0000","0000","0000","0000","0000","0000","0010","0110","1101","1101","0110","0011","0001","0000","0010","1011","0010","0000","0001","1000","0011","0000","0000","0011","0100","0100","0100","0011","0011","0010","0000","0000","0000","0000","0000","0010","1011","0010","0000","0001","0111","0110","0110","0111","0000","0000","0100","1010","0001","0000","0000","0000","0000","0000","0001","1000","0101","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0010","1010","0010","0000","0000","0001","1011","0001","0000","0000","0011","0110","0110","0111","1000","1001","1100","0101","0000","0000","0000","0000","0001","0011","1000","1111","1000","0101","0001","0000","0000","0000","0000","0000","0000","0010","0110","1100","1101","0110","0011","0001","0000","0010","1011","0010","0000","0001","1000","0011","0000","0100","1010","1011","1011","1011","1011","1011","1001","0100","0000","0000","0000","0001","0110","0111","0001","0000","0010","1011","0010","0010","1001","0010","0000","0010","1010","0100","0000","0000","0000","0000","0000","0001","1010","0011","0000","0000","0011","0101","0001","0000","0000","0000","0000","0000","0010","0101","0001","0000","0001","1010","0011","0000","0000","0001","1010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0101","1001","0000","0000","0000","0000","0001","0011","1000","1111","1000","0101","0001","0000","0000","0000","0000","0000","0000","0010","0110","1100","1101","0110","0011","0001","0000","0010","1011","0010","0000","0001","1000","0010","0000","1000","0110","0010","0010","0001","0010","0010","0101","1001","0010","0000","0000","0001","1001","0100","0000","0000","0110","1000","0010","0010","1001","0011","0000","0000","0111","1000","0001","0000","0000","0000","0000","0010","1010","0010","0000","0001","1001","1011","0011","0000","0000","0000","0000","0001","0111","1100","0011","0000","0000","1000","0101","0000","0000","0001","1010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0101","1001","0000","0000","0000","0000","0001","0011","1000","1111","1000","0101","0001","0000","0000","0000","0000","0000","0000","0010","0110","1100","1101","0110","0011","0001","0000","0010","1011","0010","0000","0001","1000","0010","0000","1001","0100","0001","0000","0000","0000","0000","0001","1001","0011","0000","0000","0100","1010","0001","0000","0000","0110","1011","1001","1001","1010","0101","0000","0000","0011","1010","0010","0000","0000","0000","0000","0011","1010","0001","0000","0010","1010","1000","0110","0000","0000","0000","0000","0010","1011","1000","0101","0000","0000","0110","0111","0000","0000","0001","1011","0000","0000","0000","0010","0011","0011","0011","0011","0011","1010","0101","0000","0000","0000","0000","0001","0011","1000","1111","1000","0101","0010","0000","0000","0000","0000","0000","0001","0010","0101","1100","1101","0110","0011","0010","0000","0010","1011","0010","0000","0001","1000","0011","0000","0111","1000","0101","0100","0010","0000","0000","0001","1000","0100","0000","0000","0111","0110","0000","0000","0000","0010","0101","0110","0110","0110","0010","0000","0000","0001","1001","0100","0000","0000","0000","0000","0110","0111","0000","0000","0011","1010","0100","1001","0001","0000","0000","0000","0100","1001","0101","0111","0000","0000","0011","1010","0001","0000","0001","1011","0001","0000","0000","1000","1010","1010","1010","1010","1010","1001","0001","0000","0000","0000","0000","0001","0011","0111","1111","1000","0101","0010","0000","0000","0000","0000","0000","0001","0010","0101","1100","1101","0110","0100","0001","0000","0010","1011","0010","0000","0001","1001","0010","0000","0010","1000","1011","1011","1001","0001","0000","0000","1001","0100","0000","0010","1010","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0110","1000","0001","0000","0000","0000","0111","0101","0000","0000","0101","0111","0011","1011","0011","0000","0000","0000","0111","0110","0011","1001","0000","0000","0010","1010","0010","0000","0001","1010","0001","0000","0000","1011","0011","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0001","0011","0111","1111","1000","0101","0010","0000","0000","0000","0000","0000","0001","0010","0101","1100","1101","0110","0011","0001","0000","0001","1011","0011","0000","0000","0111","0110","0000","0000","0001","0011","0101","1001","0001","0000","0010","1010","0010","0000","0101","1001","0000","0000","0000","0001","0001","0001","0001","0000","0001","0000","0000","0000","0000","0010","1011","0010","0000","0000","0010","1001","0011","0000","0000","0111","0101","0001","1000","0101","0000","0000","0010","1001","0011","0001","1010","0001","0000","0001","1001","0011","0000","0001","1011","0000","0000","0001","1011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0011","0111","1111","1000","0101","0010","0000","0000","0000","0000","0000","0001","0010","0101","1100","1110","0110","0011","0001","0000","0001","1001","0100","0000","0000","0010","1010","0111","0010","0010","0100","1010","0101","0000","0000","0010","1011","0010","0001","1000","0100","0000","0000","0010","1000","1000","1000","1000","1000","1000","0111","0110","0001","0000","0000","1001","0101","0001","0000","0010","1010","0010","0000","0001","1000","0011","0000","0100","1010","0110","0100","1000","1000","0001","0001","1001","0010","0000","0000","1000","0100","0000","0001","1011","0000","0000","0001","1011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0011","0111","1111","1000","0101","0010","0000","0000","0000","0000","0000","0000","0010","0101","1100","1110","0110","0100","0001","0000","0000","0101","1000","0001","0000","0000","0011","1010","1100","1011","1100","0110","0001","0000","0000","0110","1000","0001","0010","1001","0001","0000","0000","0111","1001","0111","0111","0111","0111","1000","1001","1011","0011","0000","0000","0100","1001","0010","0000","0011","1010","0001","0000","0001","1010","0001","0000","0001","0101","1010","1100","1001","0010","0000","0001","1000","0011","0000","0000","0110","0110","0000","0001","1010","0001","0000","0001","1011","0101","0011","0011","0011","0011","0010","0010","0000","0000","0000","0000","0001","0011","0111","1111","1000","0101","0010","0000","0000","0000","0000","0000","0000","0010","0101","1100","1110","0110","0100","0001","0000","0000","0001","1010","0110","0001","0000","0000","0010","0100","0100","0011","0001","0000","0000","0011","1010","0011","0000","0110","0111","0000","0000","0010","1010","0100","0001","0001","0001","0001","0000","0001","0110","0111","0000","0000","0001","1010","0011","0000","0110","1000","0000","0000","0010","1001","0001","0000","0000","0001","0010","0010","0010","0000","0000","0000","0111","0101","0000","0000","0100","1001","0001","0001","1011","0000","0000","0000","0110","1011","1011","1011","1010","1011","1011","1010","0110","0000","0000","0000","0001","0011","0111","1111","1000","0101","0010","0000","0000","0000","0000","0000","0000","0010","0101","1100","1110","0111","0100","0001","0000","0000","0000","0011","1011","0100","0001","0000","0000","0000","0000","0000","0000","0000","0010","1001","0111","0001","0001","1001","0100","0000","0000","0100","1001","0001","0000","0000","0000","0000","0000","0000","0011","1011","0010","0000","0000","0111","0100","0000","0110","0101","0000","0000","0100","1001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0110","0111","0000","0000","0010","1010","0010","0001","1010","0001","0000","0000","0000","0001","0001","0001","0010","0010","0001","0011","1011","0001","0000","0000","0001","0010","0111","1111","1000","0101","0010","0000","0000","0000","0000","0000","0000","0010","0101","1100","1110","0111","0100","0001","0000","0000","0000","0001","0101","1011","0101","0010","0001","0000","0000","0001","0010","0100","1010","1001","0010","0000","0000","1000","0110","0001","0010","1000","0110","0000","0000","0000","0000","0000","0000","0000","0010","1001","0101","0000","0001","1000","0100","0000","0110","0110","0001","0001","0111","0111","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0100","1001","0010","0000","0010","1010","0010","0001","1010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1010","0010","0000","0000","0001","0010","0111","1111","1000","0101","0010","0000","0000","0000","0000","0000","0000","0001","0101","1100","1110","0111","0100","0010","0001","0000","0000","0000","0001","0100","1010","1010","1000","1000","0111","0111","1010","1010","0111","0010","0000","0000","0000","0100","1010","1000","1010","1000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0101","1011","0111","0111","1010","0010","0000","0011","1010","1000","1000","1010","0011","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","1010","1000","0101","0111","1001","0001","0000","1001","0111","0010","0010","0010","0010","0001","0001","0001","0001","0001","0011","1011","0001","0000","0000","0001","0010","0111","1111","1000","0101","0010","0000","0000","0000","0000","0000","0000","0001","0101","1011","1110","0111","0100","0010","0001","0000","0000","0000","0000","0001","0010","0101","0111","1000","1001","1000","0101","0011","0001","0000","0000","0000","0000","0001","0100","1000","0101","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0101","1000","1001","0100","0000","0000","0001","0100","0111","0111","0100","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0100","1010","1100","1010","0011","0000","0000","0010","1011","1101","1101","1100","1101","1100","1100","1100","1100","1100","1100","0111","0000","0000","0000","0001","0010","0111","1111","1000","0101","0010","0000","0000","0000","0000","0000","0000","0001","0101","1011","1110","0111","0100","0010","0001","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0001","0001","0000","0000","0000","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0010","0001","0000","0000","0000","0000","0001","0100","0100","0100","0100","0101","0100","0100","0101","0101","0100","0000","0000","0000","0000","0001","0010","0111","1111","1000","0101","0010","0000","0000","0000","0000","0000","0000","0001","0100","1011","1110","0110","0100","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0111","1111","1000","0101","0010","0000","0000","0000","0000","0000","0000","0001","0100","1011","1110","0110","0100","0001","0001","0000","0000","0000","0000","0000","0000","0000","0010","0011","0100","0100","0011","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0111","1111","1000","0101","0010","0000","0000","0000","0000","0000","0000","0001","0100","1010","1110","0110","0100","0010","0001","0000","0000","0000","0000","0001","0100","1000","1010","1010","1010","1011","1010","1010","1001","0100","0000","0000","0000","0000","0000","0001","0111","1010","1000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1000","1001","0100","0000","0000","0000","0001","0101","1001","1000","1000","1000","1000","1000","1000","1000","1000","1000","0111","0011","0000","0000","0000","0010","0110","1000","1000","1000","1000","1000","1000","0110","0110","0100","0010","0000","0000","0000","0000","0000","0000","0000","0001","0010","0111","1111","1000","0101","0010","0000","0000","0000","0001","0001","0000","0001","0100","1010","1110","0110","0011","0001","0001","0000","0000","0000","0001","0110","1011","0111","0011","0001","0001","0000","0001","0011","0111","1100","0110","0000","0000","0000","0000","0111","1001","0101","1001","1001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1011","1000","0111","1011","0011","0000","0000","0100","1011","0110","0101","0101","0101","0101","0101","0101","0101","0101","0110","0111","1010","0001","0000","0000","0111","1010","0110","0101","0101","0110","0110","0101","0111","1000","1011","1001","0011","0001","0000","0000","0000","0000","0000","0001","0010","0111","1111","1000","0101","0010","0000","0000","0000","0000","0000","0000","0001","0100","1010","1110","0110","0011","0001","0000","0000","0000","0000","0101","1100","0011","0000","0000","0000","0000","0000","0000","0000","0000","0100","1011","0110","0000","0000","0000","1010","0010","0000","0001","1011","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0101","1001","0001","0000","0101","1000","0000","0001","1010","0101","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1001","0011","0000","0001","1001","0011","0000","0000","0000","0000","0000","0000","0000","0001","0010","1000","1011","0101","0001","0000","0000","0000","0000","0001","0010","0111","1111","1000","0101","0010","0000","0000","0000","0000","0000","0000","0001","0100","1010","1110","0110","0011","0001","0000","0000","0000","0101","1011","0011","0000","0000","0000","0001","0010","0010","0001","0000","0000","0000","0011","1010","0101","0000","0000","1010","0001","0000","0000","0111","0111","0000","0000","0000","0000","0001","0000","0000","0000","0000","1001","0100","0000","0000","0101","1001","0000","0011","1001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1010","0011","0000","0001","1001","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0101","1011","0100","0000","0000","0000","0000","0000","0010","0110","1111","1000","0101","0010","0001","0000","0000","0000","0000","0000","0001","0101","1011","1110","0110","0011","0001","0000","0000","0001","1010","0101","0000","0000","0000","0100","1010","1101","1101","1011","0101","0000","0000","0000","0101","1011","0001","0000","1000","0011","0000","0000","0011","1010","0001","0000","0000","0000","0000","0001","0000","0000","0001","1011","0001","0000","0000","1001","0101","0000","0011","1001","0001","0000","0000","0010","0011","0011","0011","0011","0011","0011","0010","0100","1011","0001","0000","0001","1010","0010","0000","0000","0011","0101","0101","0100","0011","0010","0000","0000","0001","0101","1010","0001","0000","0000","0000","0000","0010","0110","1111","1001","0110","0010","0001","0000","0000","0000","0000","0000","0001","0101","1010","1110","0110","0011","0001","0000","0000","0101","1001","0001","0000","0000","0101","1011","1000","0101","0100","0111","1011","0111","0000","0000","0000","1000","0110","0000","0101","1000","0000","0000","0001","1010","0010","0000","0000","0000","0000","0000","0000","0000","0101","1001","0000","0000","0001","1011","0001","0000","0011","1001","0001","0000","0001","1000","1011","1100","1011","1011","1011","1010","1011","1011","0101","0001","0000","0001","1010","0010","0000","0001","1001","1010","1011","1011","1011","1001","0100","0000","0000","0001","1001","0100","0000","0000","0000","0000","0010","0110","1111","1001","0110","0010","0001","0000","0000","0000","0000","0000","0001","0101","1010","1110","0110","0011","0001","0000","0000","1001","0100","0000","0000","0011","1011","0100","0000","0000","0000","0000","0011","1010","0100","0000","0000","0011","1010","0000","0001","1010","0001","0000","0000","0111","0110","0000","0000","0000","0000","0000","0000","0000","1010","0011","0000","0000","0101","1001","0000","0000","0011","1001","0001","0000","0010","1011","0100","0001","0010","0010","0010","0010","0010","0010","0001","0000","0000","0001","1010","0001","0000","0001","1001","0011","0001","0001","0011","0101","1010","0010","0000","0000","0100","1001","0000","0000","0000","0000","0010","0110","1111","1001","0110","0010","0001","0000","0000","0000","0000","0000","0001","0101","1010","1111","0110","0011","0001","0000","0001","1011","0001","0000","0000","1001","0101","0000","0000","0000","0000","0000","0000","0100","1001","0000","0000","0001","1010","0001","0000","1000","0100","0000","0000","0011","1010","0001","0000","0000","0000","0000","0000","0010","1011","0000","0000","0000","1001","0100","0000","0000","0011","1001","0001","0000","0010","1011","0010","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0001","1001","0001","0000","0000","1001","0010","0000","0000","0000","0001","1000","0100","0000","0000","0010","1011","0010","0000","0000","0000","0010","0110","1111","1001","0110","0010","0001","0000","0000","0000","0000","0000","0001","0100","1010","1111","0110","0011","0001","0000","0001","1011","0001","0000","0000","1010","0001","0000","0000","0000","0000","0000","0000","0010","1001","0000","0000","0001","1011","0001","0000","0100","1001","0000","0000","0000","1010","0011","0000","0000","0000","0000","0000","0111","0111","0000","0000","0010","1011","0001","0000","0000","0011","1000","0001","0000","0010","1011","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1010","0001","0000","0001","1001","0010","0000","0000","0000","0000","0111","0110","0000","0000","0001","1010","0010","0000","0000","0000","0010","0110","1111","1001","0110","0010","0001","0000","0000","0000","0000","0000","0001","0100","1010","1111","0110","0011","0001","0000","0001","1011","0000","0000","0001","1010","0001","0000","0000","0000","0000","0000","0000","0010","1010","0000","0000","0001","1011","0000","0000","0001","1011","0010","0000","0000","0111","0110","0000","0000","0000","0000","0001","1011","0010","0000","0000","0110","0111","0000","0000","0000","0011","1000","0001","0000","0011","1011","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1001","0010","0000","0001","1001","0010","0000","0000","0000","0000","0110","0110","0000","0000","0001","1010","0010","0000","0000","0000","0010","0110","1111","1001","0110","0010","0001","0000","0000","0000","0000","0000","0001","0100","1010","1111","0110","0011","0001","0000","0001","1100","0001","0000","0001","1011","0000","0000","0000","0000","0000","0000","0000","0001","1010","0000","0000","0001","1011","0001","0000","0000","1000","0101","0000","0000","0011","1010","0001","0000","0000","0000","0100","1010","0000","0000","0000","1010","0011","0000","0000","0000","0011","1001","0001","0000","0010","1011","0011","0011","0011","0010","0010","0010","0001","0001","0000","0000","0000","0001","1010","0001","0000","0001","1001","0010","0000","0000","0000","0010","1010","0011","0000","0000","0010","1010","0010","0000","0000","0000","0010","0110","1111","1001","0110","0010","0001","0000","0000","0000","0000","0000","0001","0100","1010","1111","0110","0011","0001","0000","0001","1011","0000","0000","0001","1011","0001","0000","0000","0000","0000","0000","0000","0001","1010","0000","0000","0001","1011","0001","0000","0000","0100","1001","0000","0000","0001","1010","0011","0000","0000","0000","0111","0110","0000","0000","0100","1010","0001","0000","0000","0000","0011","1001","0001","0000","0001","0111","1010","1010","1010","1011","1010","1010","1001","0010","0000","0000","0000","0010","1010","0001","0000","0001","1010","0101","0011","0011","0101","1001","1000","0001","0000","0000","0100","1001","0001","0000","0000","0001","0010","0110","1111","1001","0110","0010","0001","0000","0000","0000","0000","0000","0001","0100","1010","1111","0110","0011","0001","0000","0001","1011","0000","0000","0001","1011","0001","0000","0000","0000","0000","0000","0000","0010","1010","0000","0000","0001","1011","0001","0000","0000","0001","1011","0001","0000","0000","0110","0111","0000","0000","0001","1011","0010","0000","0000","0111","0110","0000","0000","0000","0000","0011","1001","0001","0000","0000","0001","0011","0011","0011","0011","0100","0011","1001","0100","0000","0000","0000","0001","1010","0010","0000","0001","1010","1100","1101","1101","1100","0111","0010","0000","0000","0001","0111","0110","0000","0000","0000","0001","0010","0110","1111","1001","0110","0010","0001","0000","0000","0000","0000","0000","0001","0100","1010","1111","0110","0011","0001","0000","0001","1011","0000","0000","0001","1011","0001","0000","0000","0000","0000","0000","0000","0010","1010","0000","0000","0001","1011","0001","0000","0000","0000","0111","0110","0000","0000","0010","1010","0001","0000","0100","1000","0000","0000","0001","1011","0010","0000","0000","0000","0000","0011","1000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0101","1000","0000","0000","0000","0010","1010","0010","0000","0000","0010","0011","0011","0010","0010","0001","0000","0000","0000","0011","1011","0010","0000","0000","0000","0000","0010","0110","1111","1001","0110","0010","0001","0000","0000","0000","0000","0000","0001","0100","1010","1111","0110","0011","0001","0000","0001","1011","0000","0000","0001","1011","0001","0000","0000","0000","0000","0000","0000","0010","1010","0000","0000","0001","1011","0001","0000","0000","0000","0010","1010","0001","0000","0000","1010","0100","0000","1000","0100","0000","0000","0100","1001","0001","0001","0001","0001","0000","0100","1001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0110","0110","0000","0000","0000","0010","1010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","1000","0111","0001","0000","0000","0000","0000","0010","0110","1111","1010","0110","0010","0001","0000","0000","0000","0000","0000","0001","0100","1010","1111","0110","0011","0001","0000","0010","1011","0000","0000","0001","1011","0001","0000","0000","0000","0000","0000","0000","0001","1010","0000","0000","0001","1011","0001","0000","0000","0000","0000","1010","0010","0000","0000","0110","1000","0001","1010","0001","0000","0000","1001","0100","0000","0000","0000","0000","0000","0100","1001","0001","0000","0001","0100","0101","0101","0101","0101","0101","0101","1010","0011","0000","0000","0000","0010","1011","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1100","0011","0000","0000","0000","0000","0000","0010","0110","1111","1010","0110","0010","0001","0000","0000","0000","0000","0000","0001","0100","1010","1111","0110","0011","0001","0000","0010","1011","0000","0000","0001","1011","0001","0000","0000","0000","0000","0000","0000","0010","1010","0000","0000","0000","1011","0001","0000","0000","0000","0000","0111","0111","0000","0000","0010","1010","0111","1000","0000","0000","0010","1011","0001","0000","0000","0000","0000","0000","0011","1001","0000","0000","0010","1010","1001","1001","1001","1001","1001","1000","0101","0001","0000","0000","0000","0010","1011","0010","0000","0000","0100","0110","0110","0110","0110","0101","0000","0000","0001","1000","0111","0000","0000","0000","0000","0000","0010","0110","1111","1010","0110","0010","0001","0000","0000","0000","0000","0000","0001","0100","1010","1111","0110","0011","0001","0000","0010","1011","0000","0000","0001","1011","0001","0000","0000","0000","0000","0000","0000","0010","1010","0000","0000","0001","1011","0001","0000","0000","0000","0000","0010","1011","0000","0000","0000","0111","1010","0010","0000","0000","0101","1000","0000","0000","0000","0000","0000","0000","0011","1000","0000","0000","0010","1011","0010","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0001","1010","0010","0000","0001","1001","1001","1001","1001","1001","1011","0011","0000","0000","0011","1010","0010","0000","0000","0000","0000","0010","0110","1111","1010","0110","0010","0001","0000","0000","0000","0000","0000","0010","0101","1010","1111","0110","0011","0001","0000","0010","1011","0000","0000","0001","1011","0001","0000","0000","0000","0000","0000","0000","0011","1010","0000","0000","0001","1011","0001","0000","0000","0000","0000","0000","1010","0010","0000","0000","0001","0010","0000","0000","0000","1001","0011","0000","0000","0000","0000","0000","0000","0011","1000","0001","0000","0010","1011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","1010","0001","0000","0001","1001","0010","0001","0001","0001","0110","1001","0001","0000","0001","1001","0010","0000","0000","0000","0001","0010","0110","1111","1010","0110","0010","0001","0000","0000","0000","0000","0000","0010","0101","1010","1111","0110","0011","0001","0000","0001","1011","0000","0000","0000","1001","0101","0000","0000","0000","0000","0000","0001","1001","0101","0000","0000","0010","1011","0001","0000","0000","0000","0000","0000","0110","1000","0000","0000","0000","0000","0000","0000","0010","1011","0000","0000","0000","0000","0000","0000","0000","0011","1000","0000","0000","0010","1011","0010","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0010","1010","0001","0000","0001","1001","0001","0000","0000","0000","0010","1011","0010","0000","0000","1001","0011","0000","0000","0001","0001","0010","0110","1111","1010","0101","0010","0001","0001","0000","0000","0000","0000","0010","0101","1010","1111","0110","0011","0001","0000","0001","1010","0010","0000","0000","0100","1011","0011","0000","0000","0000","0000","0110","1011","0001","0000","0000","0100","1010","0000","0000","0000","0000","0000","0000","0011","1010","0001","0000","0000","0000","0000","0000","0111","0111","0000","0000","0000","0000","0000","0000","0000","0100","1001","0000","0000","0010","1011","0010","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0010","1010","0001","0000","0001","1001","0001","0000","0000","0000","0001","1010","0010","0000","0001","1000","0011","0000","0000","0001","0001","0010","0110","1111","1010","0101","0010","0001","0001","0000","0000","0000","0000","0010","0101","1001","1111","0110","0011","0010","0001","0001","0110","0111","0000","0000","0000","0110","1011","0111","0101","0110","1000","1010","0011","0000","0000","0000","1001","0110","0000","0000","0000","0000","0000","0001","0000","1001","0011","0000","0000","0000","0000","0001","1011","0011","0000","0000","0000","0000","0000","0000","0000","0011","1000","0001","0000","0010","1011","0011","0010","0011","0011","0010","0010","0010","0010","0001","0000","0000","0010","1010","0001","0000","0001","1001","0010","0000","0000","0000","0001","1010","0010","0000","0001","1001","0100","0000","0000","0000","0001","0010","0110","1111","1010","0101","0010","0001","0000","0000","0000","0000","0000","0010","0101","1001","1111","0110","0011","0001","0001","0001","0010","1011","0011","0000","0000","0000","0100","0111","1001","1001","0110","0001","0000","0000","0000","0110","1010","0001","0000","0000","0000","0000","0001","0000","0000","0101","0111","0000","0000","0001","0000","0100","1010","0000","0000","0000","0000","0000","0000","0000","0000","0100","1001","0000","0000","0001","1000","1100","1100","1100","1011","1100","1011","1010","1001","0011","0000","0000","0010","1010","0000","0000","0001","1010","0010","0000","0000","0000","0001","1010","0010","0000","0000","1000","0100","0000","0000","0000","0000","0010","0110","1111","1010","0110","0010","0001","0000","0000","0000","0000","0000","0010","0101","1001","1111","0101","0010","0001","0001","0001","0000","0101","1011","0011","0000","0000","0000","0000","0001","0001","0000","0000","0000","0000","0100","1100","0100","0000","0001","0000","0000","0000","0000","0000","0000","0010","1011","0000","0000","0001","0000","1000","0110","0000","0000","0000","0001","0000","0000","0000","0000","0100","1000","0001","0000","0000","0001","0011","0011","0100","0101","0100","0101","0101","0110","1010","0001","0000","0010","1010","0001","0000","0010","1001","0001","0000","0000","0000","0001","1001","0011","0000","0001","0111","0101","0000","0000","0000","0000","0010","0101","1111","1011","0110","0011","0001","0000","0000","0000","0000","0000","0010","0101","1001","1111","0101","0011","0001","0001","0001","0000","0000","0101","1010","0101","0001","0000","0000","0000","0000","0000","0000","0001","0110","1010","0101","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","1001","0101","0000","0000","0010","1011","0010","0000","0000","0000","0000","0000","0000","0000","0000","0100","1001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1010","0010","0000","0010","1011","0001","0000","0001","1010","0010","0000","0000","0000","0001","1001","0010","0000","0000","0111","0101","0000","0000","0000","0000","0010","0110","1111","1011","0110","0011","0001","0000","0000","0000","0000","0001","0010","0101","1001","1111","0110","0011","0001","0001","0000","0000","0000","0000","0100","1100","1000","0011","0001","0000","0000","0001","0011","1001","1100","0100","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0101","1010","0010","0010","0111","1000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0011","1010","0010","0001","0000","0001","0000","0000","0000","0000","0000","0001","0001","0010","1011","0011","0000","0010","1011","0010","0001","0010","1010","0010","0000","0000","0000","0001","1001","0100","0001","0001","1000","0100","0000","0000","0000","0001","0010","0110","1111","1011","0110","0010","0001","0000","0000","0000","0000","0001","0010","0101","1001","1111","0110","0011","0010","0001","0000","0000","0000","0000","0000","0011","1001","1011","1001","1001","1001","1010","1011","1000","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","1001","1011","1010","1010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0111","1010","0111","0111","0111","0110","0110","0111","0110","0111","0111","0111","1000","1000","0001","0000","0001","1010","1000","0110","1001","1000","0001","0000","0000","0000","0000","0110","1001","0110","0110","1010","0001","0000","0000","0000","0001","0011","0110","1111","1011","0110","0010","0001","0000","0000","0000","0000","0001","0010","0100","1001","1111","0111","0100","0010","0001","0001","0000","0000","0000","0000","0000","0000","0010","0011","0100","0100","0100","0010","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0101","0110","0110","0110","0110","0110","0110","0110","0110","0111","0110","0101","0010","0000","0000","0000","0011","0110","0111","0110","0010","0000","0000","0000","0000","0000","0010","0110","1000","0111","0011","0000","0000","0000","0000","0001","0010","0110","1110","1011","0110","0010","0001","0000","0000","0000","0000","0000","0001","0100","1000","1111","1000","0110","0100","0010","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0010","0001","0001","0000","0000","0000","0000","0000","0010","0010","0110","1111","1011","0110","0010","0001","0000","0000","0000","0000","0000","0001","0011","0110","1111","1011","0111","0110","0101","0100","0010","0001","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0001","0001","0010","0001","0010","0001","0010","0001","0010","0010","0001","0001","0000","0000","0000","0001","0001","0001","0001","0000","0000","0000","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0010","0010","0011","0110","1111","1010","0101","0010","0000","0000","0000","0000","0000","0000","0000","0001","0100","1011","1111","1010","1000","0110","0110","0100","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0010","0011","0011","0011","0100","0011","0011","0100","0011","0011","0010","0001","0001","0000","0001","0011","0011","0011","0010","0001","0001","0001","0001","0010","0010","0010","0011","0011","0011","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0010","0011","0010","0010","0010","0010","0010","0010","0001","0001","0010","0001","0001","0000","0001","0001","0001","0001","0001","0001","0000","0000","0000","0001","0001","0010","0100","0101","1000","1111","1000","0101","0010","0000","0000","0000","0000","0000","0000","0000","0001","0011","0110","1101","1111","1101","1011","1001","0111","0101","0010","0010","0011","0101","0101","0100","0010","0010","0010","0011","0101","0111","0111","0111","0111","0111","0110","0111","0111","0110","0111","0101","0010","0010","0001","0011","0101","0110","0110","0101","0011","0010","0010","0011","0101","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0110","0101","0101","0101","0100","0100","0100","0011","0010","0001","0010","0011","0100","0011","0011","0001","0000","0000","0001","0010","0100","0100","0111","1000","1101","1101","0111","0011","0001","0000","0000","0000","0000","0000","0000","0000","0001","0010","0011","0110","1011","1110","1111","1111","1111","1001","0100","0011","0110","1011","1110","1011","0110","0011","0011","0110","1100","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1011","0100","0011","0011","0101","1010","1110","1101","1000","0100","0011","0011","0101","1010","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1100","1100","1100","1100","1100","1100","1100","1100","1100","1100","1011","1011","1011","1010","1010","0110","0011","0010","0100","0111","1001","1000","0100","0011","0000","0000","0010","0100","1000","1010","1011","1111","1111","1000","0101","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0011","0100","0101","0111","1001","1010","1110","1110","0110","0101","1000","1111","1101","1111","1010","0101","0110","1001","1111","1101","1101","1101","1101","1101","1101","1101","1101","1101","1101","1111","1000","0100","0100","1010","1111","1110","1111","1111","1000","0100","0101","1001","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1111","1010","0100","0011","0111","1111","1111","1111","1001","0100","0010","0010","0100","1000","1111","1111","1111","1110","1001","0110","0101","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0011","0011","0110","0111","1011","1111","0111","0110","1011","1111","1001","1100","1110","0111","0111","1011","1111","1000","1000","1000","1000","0111","0111","1000","1000","1000","1000","1111","1000","0101","0111","1101","1100","1000","1001","1111","1010","0110","0101","1100","1101","1001","1000","1000","1000","0111","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1000","1001","1100","1111","0110","0101","1011","1110","1001","1100","1110","0101","0011","0010","0101","1100","1101","1001","1000","1000","0110","0101","0100","0010","0001","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0001","0001","0011","0101","1010","1111","0111","0110","1011","1111","1000","1011","1111","1000","1000","1011","1111","0111","0101","0100","0100","0100","0100","0100","0100","0101","1000","1111","1001","0110","0110","1111","1010","0111","0111","1110","1011","0110","0111","1100","1101","1000","0110","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0101","0111","1010","1111","1000","0111","1100","1101","1000","1010","1111","0110","0011","0010","0101","1101","1100","1000","0110","0100","0100","0011","0010","0001","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0101","1010","1111","0111","0110","1100","1111","1000","1001","1111","1001","1001","1101","1110","0110","0100","0010","0010","0010","0010","0010","0011","0100","0111","1111","1010","0110","0110","1110","1010","0111","0111","1110","1011","0111","0111","1101","1101","0111","0101","0100","0011","0010","0011","0011","0011","0011","0011","0011","0011","0011","0011","0100","0100","0100","0100","0011","0011","0011","0011","0100","0101","0101","1001","1111","1000","1000","1110","1101","1000","1010","1111","0110","0011","0010","0110","1101","1100","0111","0100","0011","0010","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0101","1010","1111","0111","0111","1011","1110","1000","1000","1111","1111","1111","1111","1011","0101","0011","0001","0001","0001","0001","0001","0010","0100","0111","1111","1010","0110","0110","1111","1011","0111","0111","1110","1100","0111","0111","1101","1100","0110","0100","0010","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0001","0010","0001","0001","0001","0001","0001","0001","0010","0010","0011","0100","1000","1111","1001","1001","1111","1100","0111","1001","1111","0111","0100","0011","0110","1101","1100","0110","0011","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0101","1010","1111","1000","0110","1100","1110","0111","0110","1000","1011","1100","1010","0110","0011","0010","0001","0000","0000","0001","0001","0001","0011","0111","1111","1001","0110","0110","1111","1011","0111","0111","1101","1100","0111","0111","1101","1011","0101","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0000","0000","0001","0000","0001","0001","0001","0010","0100","0111","1111","1111","1111","1111","1001","0111","1001","1111","0111","0100","0011","0110","1110","1011","0110","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0100","1010","1110","1000","0111","1100","1111","0111","0101","0101","0100","0101","0100","0011","0010","0001","0000","0000","0000","0000","0001","0001","0011","0110","1111","1001","0110","0111","1111","1011","0111","0111","1100","1101","1000","1000","1110","1011","0110","0011","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0000","0000","0000","0000","0000","0000","0001","0010","0011","0101","1001","1110","1111","1010","0111","0110","1000","1111","0111","0100","0100","0111","1110","1011","0110","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0100","1001","1111","1000","1000","1101","1110","0110","0011","0011","0010","0010","0001","0001","0001","0000","0000","0000","0000","0000","0001","0001","0011","0111","1111","1001","0110","0111","1111","1010","0111","0110","1001","1111","1111","1110","1111","1001","0101","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0000","0000","0000","0000","0000","0000","0001","0001","0011","0100","0101","0111","0111","0110","0110","0110","1000","1111","0111","0100","0100","0111","1110","1011","0110","0010","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0001","0011","1000","1111","1011","1010","1111","1011","0101","0011","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0011","0111","1111","1001","0110","0111","1111","1010","0110","0100","0110","1010","1110","1110","1010","0110","0100","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0011","0100","0100","0101","0100","0100","0101","1000","1111","0110","0100","0100","0111","1110","1011","0110","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0101","1011","1111","1111","1110","0111","0100","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0011","0110","1111","1001","0111","0111","1111","1010","0101","0011","0100","0110","0111","0111","0110","0100","0011","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0010","0011","0011","0010","0011","0101","1000","1111","0111","0100","0100","0111","1110","1011","0110","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0011","0101","0111","1000","0110","0100","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0110","1111","1001","0111","1000","1111","1010","0101","0010","0010","0011","0100","0100","0100","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0101","0111","1111","0111","0101","0101","0111","1110","1011","0110","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0011","0100","0100","0011","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0101","1111","1011","1001","1001","1111","1001","0100","0001","0001","0010","0011","0010","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0100","1000","1111","1001","0110","0110","1000","1111","1001","0101","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0010","0010","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0100","1010","1111","1111","1111","1111","0111","0011","0001","0000","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0011","0110","1101","1110","1010","1001","1101","1111","0111","0100","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0010","0110","1010","1110","1101","1000","0101","0010","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0100","1000","1111","1111","1111","1111","1000","0101","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0011","0101","0110","0110","0101","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0000","0000","0000","0000","0000","0000","0001","0001","0000","0000","0000","0001","0010","0101","0111","1001","1001","0111","0101","0011","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0010","0011","0011","0010","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0011","0100","0101","0100","0100","0010","0010","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0010","0011","0010","0010","0001","0001","0001","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001","0001","0001","0001","0001","0000","0000","0000","0001","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000");

begin

process(clk) begin
    if(rising_edge(clk)) then
        if(clk_counter < 1) then
            clk_counter <= clk_counter + 1;
        else
            clk_counter <= 0;
            sub_clk <= not sub_clk;
        end if;
    end if;
end process;

process(sub_clk) begin
    if(rising_edge(sub_clk)) then
        --Displaying The Boardrs.
        if(((V_counter >= 0 and V_counter < 10) or (V_counter >= 470 and V_counter < 480)) or ((H_counter >= 0 and H_counter < 10) or (H_counter >= 630 and H_counter < 640))) then
            R_out <= "0000";
            G_out <= "1001";
            B_out <= "1111";
        --Displaying The Left Player.
        elsif((V_counter >= (180 + left_move) and V_counter < (300 + left_move)) and (H_counter >= 20 and H_counter < 30)) then
            R_out <= "0111";
            G_out <= "0000";
            B_out <= "0111";
        --Displaying The Right Player.
        elsif((V_counter >= (180 + right_move) and V_counter < (300 + right_move)) and (H_counter >= 610 and H_counter < 620)) then
            R_out <= "0111";
            G_out <= "0000";
            B_out <= "0111";
        --Displaying The Ball.
        elsif((V_counter >= (235 + (V_ball_move / 10)) and V_counter < (245 + (V_ball_move / 10))) and (H_counter >= (315 + (H_ball_move / 10)) and H_counter < (325 + (H_ball_move / 10)))) then
            R_out <= "0111";
            G_out <= "0000";
            B_out <= "0000";
        else
            R_out <= (others => '0');
            G_out <= (others => '0');
            B_out <= (others => '0');
        end if;
        --Ending The Game.
        if(end_game) then
            --Displaying The Image.
            if((V_counter >= 190 and V_counter < 290) and (H_counter >= 270 and H_counter < 370)) then
                R_out <= image_R(image_counter);
                G_out <= image_G(image_counter);
                B_out <= image_B(image_counter);
                if(image_counter < 9999) then
                    image_counter <= image_counter + 1;
                else
                    image_counter <= 0;
                end if;
            --Displaying The Boardrs.
            elsif(((V_counter >= 0 and V_counter < 10) or (V_counter >= 470 and V_counter < 480)) or ((H_counter >= 0 and H_counter < 10) or (H_counter >= 630 and H_counter < 640))) then
                R_out <= "0000";
                G_out <= "1001";
                B_out <= "1111";
            else
                R_out <= (others => '0');
                G_out <= (others => '0');
                B_out <= (others => '0');
            end if;
            if(reset = '1') then
                H_counter <= 0;
                V_counter <= 0;
                image_counter <= 0;
                V_ball_move <= 0;
                H_ball_move <= 0;
                left_move <= 0;
                right_move <= 0;
                ball_down <= true;
                ball_right <= true;
                end_game <= false;
            end if;
        end if;
        -- Updating the Scanline and the Frame.
        if(H_counter < 800) then
            H_counter <= H_counter + 1;
            if(H_counter >= 656 and H_counter < 752) then
                H_sync <= '0';
            else
                H_sync <= '1';
            end if;
        else
            V_counter <= V_counter + 1;
            H_counter <= 0;
        end if;
        if(V_counter < 525) then
            if(V_counter >= 490 and V_counter < 492) then
                V_sync <= '0';
            else
                V_sync <= '1';
            end if;
        else
            V_counter <= 0;
            --control the movement of the left player.
            if(left_player = '0') then
                if(left_move < 170) then
                    left_move <= left_move + 5;
                else
                    left_move <= left_move;
                end if;
            else
                if(left_move > -170) then
                    left_move <= left_move - 5;
                else
                    left_move <= left_move;
                end if;
            end if;
            --control the movement of the right player.
            if(right_player = '0') then
                if(right_move < 170) then
                    right_move <= right_move + 5;
                else
                    right_move <= right_move;
                end if;
            else
                if(right_move > -170) then
                    right_move <= right_move - 5;
                else
                    right_move <= right_move;
                end if;
            end if;
            --control the movement of the ball.
            if(ball_down) then
                if(V_ball_move < 2250) then
                    V_ball_move <= V_ball_move + 25;
                else
                    V_ball_move <= V_ball_move - 25;
                    ball_down <= false;
                end if;
            else
                if(V_ball_move > -2250) then
                    V_ball_move <= V_ball_move - 25;
                else
                    V_ball_move <= V_ball_move + 25;
                    ball_down <= true;
                end if;
            end if;
            if(ball_right) then
                if((H_ball_move = 2850) and ((V_ball_move >= (right_move * 10) - 550 and V_ball_move < (right_move * 10) + 650) or (V_ball_move > (right_move * 10) - 650 and V_ball_move < (right_move * 10) + 550))) then
                    H_ball_move <= H_ball_move - 25;
                    ball_right <= false;
                elsif(H_ball_move < 3050) then
                    H_ball_move <= H_ball_move + 25;
                else
                    end_game <= true;
                    H_ball_move <= H_ball_move;
                end if;
            else
                if((H_ball_move = -2850) and ((V_ball_move >= (left_move * 10) - 550 and V_ball_move < (left_move * 10) + 650) or (V_ball_move > (left_move * 10) - 650 and V_ball_move < (left_move * 10) + 550))) then
                    H_ball_move <= H_ball_move + 25;
                    ball_right <= true;
                elsif(H_ball_move > -3050) then
                    H_ball_move <= H_ball_move - 25;
                else
                    end_game <= true;
                    H_ball_move <= H_ball_move;
                end if;
            end if;
        end if;
    end if;
end process;

end Behavioral;